  ADDER - 4 BIT ALL-74HC00-GATE BINARY ADDER WITH BIDIRECTIONAL BRIDGES
  * behavioral gate description
  * Automatic A/D insertion using bi-directional bridges

* Override the default bridges and force use of the bidi_bridge.

.control
pre_set auto_bridge_d_out =
+ ( ".model auto_bridge bidi_bridge(out_high=%g in_low='%g/2' in_high='%g/2' )"
+   "auto_bridge%d [ %s ] [ %s ] null auto_bridge" 1000 )
pre_set auto_bridge_d_in = ( $auto_bridge_d_out )
.endc

*** SUBCIRCUIT DEFINITIONS
.include 74HCng_auto.lib
.param vcc=3 tripdt=6n

.include ../adder_common.inc

.END
