VDMOS p channel output

m1 d g s b p1
.model p1 vdmosp vto=-1.2 is=10n kp=2 bv=-12 rb=1k
*d1 d s dmod
*.model dmod d  is=10n rs=0.1

vd d 0 -5
vg g 0 -5
vs s 0 0
vb b 0 0

.dc vd -15 1 0.1 vg 0 -5 -1

.control
run
plot vs#branch
.endc

.end
