* NGspice simuliert CJ bezüglich T falsch. CJ nimmt mit steigenden T ab.
.OPTION  GMIN=1E-14 tnom=27
.PROBE

.temp 127
.AC dec 100 100 1000k
VD1 In 0 Ac=1
RL in out 100k
Q1 out 0 0 0 NX

.MODEL NX NPN (IS=1.09e-16 NF=1.002 BF=135 VAF=70 IKF=1.2m ISE=5e-18 NE=1.25 CTS=100m
+ NR=1 BR=31 IKR=5u VAR=4 ISC=3e-16 NC=1.3
+ RC=1 RE=10 RB=920 RBM=305 IRB=20U
+ CJC=10F MJC=0.451 VJC=0.306
+ CJE=10F MJE=0.9 VJE=1.57
+ CJS=10p MJS=0.561 VJS=0.844
+ TR=2p TF=33.76p XTF=6.593 VTF=1.974 ITF=0.0002479 PTF=35
+ XTI=6.6 XTB=1.9 TIKF1=-4m AF=1.328 KF=29.39f)
