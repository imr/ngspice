Colpitt's Oscillator Circuit

r1 1 0 1
q1 2 1 3 qmod area = 100p
vcc 4 0 5 
rl 4 2 750
c1 2 3 500p
c2 4 3 4500p
l1 4 2 5uH
re 3 6 4.65k
vee 6 0 dc -15 pwl 0 -15 1e-9 -10 

.tran 30n 12u
.print tran v(2)

.model qmod nbjt level=1
+ x.mesh node=1  loc=0.0
+ x.mesh node=61 loc=3.0
+ region num=1 material=1
+ material num=1 silicon nbgnn=1e17 nbgnp=1e17
+ mobility material=1 concmod=sg fieldmod=sg
+ mobility material=1 elec major
+ mobility material=1 elec minor
+ mobility material=1 hole major
+ mobility material=1 hole minor
+ doping unif n.type conc=1e17 x.l=0.0 x.h=1.0
+ doping unif p.type conc=1e16 x.l=0.0 x.h=1.5
+ doping unif n.type conc=1e15 x.l=0.0 x.h=3.0
+ models bgnw srh conctau auger concmob fieldmob
+ options base.length=1.0 base.depth=1.25

.options acct bypass=1
.end
