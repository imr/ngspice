***  For BSIM3V3.1 general purpose check (Id-Vd) for Pmosfet ***
******************************************

*** circuit description ***
m1 2 1 0 0 p1 L=0.35u W=10.0u
vgs 1 0 -3.5
vds 2 0 -3.5

.options noacct
.dc vds 0 -3.5 -0.05 vgs 0 -3.5 -0.5


.print dc v(1) i(vds)


.include modelcard.pmos 
.end


