DIODE REVERSE RECOVERY

VPP 1 0 0.0V (PULSE 1.0V -1.0V 1NS 1PS 1PS 20NS 40NS)
VNN 2 0 0.0V
RS  1 3 1.0
LS  3 4 0.5UH
DT  4 2 M_PIN AREA=1

.MODEL M_PIN NUMD LEVEL=2
+ OPTIONS DEFW=100U
+ X.MESH N=1 L=0.0
+ X.MESH N=2 L=0.2
+ X.MESH N=4 L=0.4
+ X.MESH N=8 L=0.6
+ X.MESH N=13 L=1.0
+
+ Y.MESH N=1 L=0.0
+ Y.MESH N=9 L=4.0
+ Y.MESH N=24 L=10.0
+ Y.MESH N=29 L=15.0
+ Y.MESH N=34 L=20.0
+
+ DOMAIN NUM=1 MATERIAL=1
+ MATERIAL NUM=1 SILICON TN=20NS TP=20NS
+
+ ELECTRODE NUM=1 X.L=0.6 X.H=1.0 Y.L=0.0 Y.H=0.0
+ ELECTRODE NUM=2 X.L=-0.1 X.H=1.0 Y.L=20.0 Y.H=20.0
+
+ DOPING GAUSS P.TYPE CONC=1.0E19 CHAR.LEN=1.076 X.L=0.75 X.H=1.1 Y.H=0.0
+ + LAT.ROTATE RATIO=0.1
+ DOPING UNIF  N.TYPE CONC=1.0E14
+ DOPING GAUSS N.TYPE CONC=1.0E19 CHAR.LEN=1.614 X.L=-0.1 X.H=1.1 Y.L=20.0
+
+ MODELS BGN SRH AUGER CONCTAU CONCMOB FIELDMOB

.OPTION ACCT BYPASS=1
.TRAN 0.1NS 10NS
.PRINT TRAN V(3) I(VIN)

.END
