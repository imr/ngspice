regression test temper-1.cir, 'temper' in a model parameter

* check inp_evaluate_temper() processing

.model dplain d is='temper+1000'

D1  1 0  dplain

.control

let success_count = 0

op

let val = @dplain[is]
let gold = 1000 + 27.0

let err = abs(val/gold - 1)

echo "Note: err =" $&err

if err > 1e-12
  echo "ERROR: test failed"
else
  echo "INFO: success"
  let success_count = success_count + 1
end

if success_count ne 1
  quit 1
else
  quit 0
end

.endc

.end
