BiCMOS Pulldown Circuit

VSS 2 0 0v

VIN 3 2 0v (PULSE 0.0v 4.2v 0ns 1ns 1ns 9ns 20ns)

M1  8 3 5 11 M_NMOS_1 W=4u L=1u
VD  4 8 0v
VBK 11 2 0v

Q1  10 7 9   M_NPN AREA=8
VC  4 10 0v
VB  5 7 0v
VE  9 2 0v

CL  4 6 1pF
VL  6 2 0v

.IC V(10)=5.0v V(7)=0.0v 
.TRAN 0.1ns 5ns 0ns 0.1ns
.PLOT TRAN I(VIN)

.include bicmos.lib

.OPTIONS ACCT BYPASS=1
.END
