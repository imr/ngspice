MOS CHARGE PUMP

VIN 4 0 DC 0V PULSE 0 5 15NS 5NS 5NS 50NS 100NS
VDD 5 6 DC 0V PULSE 0 5 25NS 5NS 5NS 50NS 100NS
VBB 0 7 DC 0V PULSE 0 5  0NS 5NS 5NS 50NS 100NS
RD 6 2 10K
M1 5 4 3 7 MMOD W=100UM
VS 3 2 0
VC 2 1 0
C2 1 0 10PF

.IC V(3)=1.0
.TRAN 2NS 200NS
.OPTIONS ACCT BYPASS=1
.PRINT TRAN V(1) V(2)

.MODEL MMOD NUMOS
+ X.MESH N=1 L=0
+ X.MESH N=3 L=0.4
+ X.MESH N=7 L=0.6
+ X.MESH N=15 L=1.4
+ X.MESH N=19 L=1.6
+ X.MESH N=21 L=2.0
+
+ Y.MESH N=1 L=0
+ Y.MESH N=4 L=0.015
+ Y.MESH N=8 L=0.05
+ Y.MESH N=12 L=0.25
+ Y.MESH N=14 L=0.35
+ Y.MESH N=17 L=0.5
+ Y.MESH N=21 L=1.0
+
+ REGION NUM=1 MATERIAL=1 Y.L=0.015
+ MATERIAL NUM=1 SILICON
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+
+ REGION NUM=2 MATERIAL=2 Y.H=0.015 X.L=0.5 X.H=1.5
+ MATERIAL NUM=2 OXIDE
+
+ ELEC NUM=1 IX.L=18 IX.H=21   IY.L=4  IY.H=4
+ ELEC NUM=2 IX.L=5  IX.H=17   IY.L=1  IY.H=1
+ ELEC NUM=3 IX.L=1  IX.H=4    IY.L=4  IY.H=4
+ ELEC NUM=4 IX.L=1  IX.H=21   IY.L=21 IY.H=21
+
+ DOPING UNIF N.TYPE CONC=1E18   X.L=0.0 X.H=0.5 Y.L=0.015 Y.H=0.25
+ DOPING UNIF N.TYPE CONC=1E18   X.L=1.5 X.H=2.0 Y.L=0.015 Y.H=0.25
+ DOPING UNIF P.TYPE CONC=1E15   X.L=0.0 X.H=2.0 Y.L=0.015 Y.H=1.0
+ DOPING UNIF P.TYPE CONC=1.3E17 X.L=0.5 X.H=1.5 Y.L=0.015 Y.H=0.05
+
+ MODELS CONCMOB FIELDMOB
+ METHOD ONEC

.END
