test pz
iin	1	0	ac
r1	1	0	1Ohms
l1	1	0	0.05H

gm2	2	0	1 0 1
r2	2	0	1Ohms
l2	2	0	0.05H

gm3	3	0	2 0 1
r3	3	0	1Ohms
l3	3	0	0.05H

*gm4	4	0	3 0 1
*r4	4	0	1Ohms
*l4	4	0	0.05H

*gm5	5	0	4 0 1
*r5	5	0	10Ohms
*l5	5	0	0.66mH

.pz	1 0	3 0	cur pol
.print pz all
.end
