* test inductor branch current, tran, without feedback
*  (exec-spice "ngspice %s" t)

V1   in 0   SINE(0 1 1)

L1   in N3  0.21 m = 3
Vm1  N3 N5  0
R2   N5 0   1.0

B1   out 0  V = I(L1)

.control

* insertion of nodes and branches has to be checked for correct "unsetup"
* I saw a failing tran after an op, whilst tran alone worked

op
rusage totiter

tran 1ms 1.0
rusage totiter

* golden answer, derived with "maxima"
let R = 1
let L = 0.21 / 3
let tau = L / R
let omega = 2 * pi
let ot = omega * tau
let gold = (sin(time*omega) - ot*cos(time*omega) + ot*exp(-time/tau)) / (1+ot*ot)/R

let err = vecmax(abs(v(out) - gold))
echo "INFO: err =" $&err

if err > 6e-6
  echo "ERROR: test failed"
  quit 1
else
  echo "INFO: success"
end

if 1
  plot v(out) i(Vm1)*0.99 v(N5)*0.98 gold*0.97
  plot v(out)-gold
else
  quit 0
end

.endc

.end
