** NMOSFET: Benchmarking Implementation of BSIM4 by Jane Xi 05/09/2003.

** Circuit Description **
m1 2 1  0 3 n1 L=0.09u W=10.0u rgeoMod=1
vgs 1 0 1.2 
vbs 3 0 0 
vds 2 0 0.1

.dc vgs -0.6 1.2 0.02 vbs 0.0 -1.2 -0.3

.options noacct

.print dc v(2) i(vds)

.include  modelcard.nmos
.end
