Example circuit to read a Touchstone-format parameter file.

* This file contains an an analog filter circuit; SP and AC analyses are run
* and the S-parameters are saved in a file.  It also contains a behavioural
* circuit that reproduces the original from its saved S-parameters.
* Results from the two versions are plotted together for comparison.
* The behavioural circuit also illustrates the use of a string-valued
* sub-circuit parameter to pass a file name.

* Derived from: Qucs 1.0.2 C:/Users/Tom Hajjar/.qucs - S/S-parameter_files_ngspice_prj/137MHz_BPF.sch

* Original circuit for SP analysis

VP2 _net0 0 dc 0 ac 0.316228 SIN(0 0.316228 1G) portnum 2 z0 50
VP1 _net1 0 dc 0 ac 0.316228 SIN(0 0.316228 1G) portnum 1 z0 50
C1 _net2 _net1  4.7P 
C5 _net3 _net0  4.7P 
C3 _net3 _net2  1P 
C4 _net3 0  15P 
C2 0 _net2  15P 
L2 0 _net3  66N 
L1 0 _net2  66N 

.csparam Rbase=50 ; This is required by "wrs2p", below.

* A version derived from extracted s-parameters, with option for subcircuit.

VP3 net1 0 dc 0 ac 0.316228 ; Same as VP1 but that must not be loaded.
ri net1 sin 50
.param in_file="137MHz_BPF.s2p"
X1 sin sout 0 s2p_generic touchstone=in_file
ro sout 0 50

* Control section, run simulations.

.control
* Run an SP analysis, derive group delay and write a Touchstone file

SP LIN 71 107MEG 167MEG
let Group_Delay = -1*deriv(cph(S_2_1))/(2*pi)
wrs2p  new_137MHz_BPF.s2p

* Now run AC analysis

alter vp2 ac = 0
AC LIN 71 107MEG 167MEG
set xbrushwidth=2
plot group_delay(_net0) sp1.Group_Delay group_delay(sout)
plot db(_net0) cph(_net0) db(sout) cph(sout)
.endc

* Subcircuit for SP behavioral device

.SUBCKT s2p_generic  1 2 3 touchstone={touchstone}
* Pin 3 is the reference plane (usually it should be connected to GND)
* HZ S RI R 50
* Z1 = 50 Z2 = 50
R1N 1 100 -5.000000e+01
R1P 100 101 100.000000
R2N 2 200 -5.000000e+01
R2P 200 201 100.000000

* S11 FREQ R_I
 A0101 %vd 100 3 %vd 101 102 m_a0101
 .model m_a0101 xfer file=touchstone span=9

* S12 FREQ R_I
 A0102 %vd 200 3 %vd 102 3 m_a0102
 .model m_a0102 xfer file=touchstone span=9 offset=3

* S21 FREQ R_I
 A0201 %vd 100 3 %vd 201 202 m_a0201
 .model m_a0201 xfer file=touchstone span=9 offset=5

* S22 FREQ R_I
 A0202 %vd 200 3 %vd 202 3 m_a0202
 .model m_a0202 xfer file=touchstone span=9 offset=7

.ENDS

.END
