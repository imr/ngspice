NMOS Enhancement-Load Bootstrap Inverter

Vdd 1 0 5.0v
Vss 2 0 0.0v

Vin 5 0 0.0v PWL (0.0ns 5.0v) (1ns 0.0v) (10ns 0.0v) (11ns 5.0v)
+ (20ns 5.0v) (21ns 0.0v) (30ns 0.0v) (31ns 5.0v)
M1  1 1 3 2 M_NMOS w=5u
M2  1 3 4 4 M_NMOS w=5u
M3  4 5 2 2 M_NMOS w=5u
CL  4 0 0.1pf
CB  3 4 0.1pf

.model M_NMOS numos
+ x.mesh l=0.0 n=1
+ x.mesh l=0.6 n=4
+ x.mesh l=0.7 n=5
+ x.mesh l=1.0 n=7
+ x.mesh l=1.2 n=11
+ x.mesh l=3.2 n=21
+ x.mesh l=3.4 n=25
+ x.mesh l=3.7 n=27
+ x.mesh l=3.8 n=28
+ x.mesh l=4.4 n=31
+
+ y.mesh l=-.05 n=1
+ y.mesh l=0.0  n=5
+ y.mesh l=.05  n=9
+ y.mesh l=0.3  n=14
+ y.mesh l=2.0  n=19
+
+ region num=1 material=1 y.l=0.0
+ material num=1 silicon
+ mobility material=1 concmod=sg fieldmod=sg
+ mobility material=1 init elec major
+ mobility material=1 init elec minor
+ mobility material=1 init hole major
+ mobility material=1 init hole minor
+
+ region num=2 material=2 y.h=0.0 x.l=0.7 x.h=3.7
+ material num=2 oxide
+
+ elec num=1 x.l=3.8 x.h=4.4	y.l=0.0 y.h=0.0
+ elec num=2 x.l=0.7 x.h=3.7	iy.l=1  iy.h=1
+ elec num=3 x.l=0.0 x.h=0.6	y.l=0.0 y.h=0.0
+ elec num=4 x.l=0.0 x.h=4.4	y.l=2.0 y.h=2.0
+
+ doping unif p.type conc=2.5e16 x.l=0.0 x.h=4.4  y.l=0.0 y.h=2.0
+ doping unif p.type conc=1e16   x.l=0.0 x.h=4.4  y.l=0.0 y.h=0.05
+ doping unif n.type conc=1e20   x.l=0.0 x.h=1.1  y.l=0.0 y.h=0.2
+ doping unif n.type conc=1e20   x.l=3.3 x.h=4.4  y.l=0.0 y.h=0.2
+
+ models concmob fieldmob
+ method ac=direct onec

.tran 0.2ns 40ns
.print v(4)
.options acct bypass=1 method=gear
.end
