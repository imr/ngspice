SWITCHED CURRENT CELL - CLOCK FEEDTHROUGH

VDD 1 0 5.0V
VSS 2 0 0.0V

IIN 13 0 0.0
VIN 13 3 0.0
VL  4 0 2.5V
VCK 6 0 5.0V PULSE 5.0V 0.0V 5.0NS 5NS 5NS 20NS 50NS

M1   3  3  2  2 M_NMOS_5 W=5U L=5U
M2   4  5  2  2 M_NMOS_5 W=10U L=5U
M3  23 26 25 22 M_NMOS_5 W=5U L=5U
RLK1 3 0 100G
RLK2 5 0 100G
VD  3 23 0.0V
VG  6 26 0.0V
VS  5 25 0.0V
VB  2 22 0.0V

M4  7 7 1 1 M_PMOS_IDEAL  W=100U L=1U
M5  3 7 1 1 M_PMOS_IDEAL  W=100U L=1U
M6  4 7 1 1 M_PMOS_IDEAL  W=200U L=1U
IREF 7 0 50UA 

****** MODELS ******
.MODEL M_PMOS_IDEAL PMOS VTO=-1.0V KP=100U

.INCLUDE BICMOS.LIB

.TRAN 0.1NS 50NS

.OPTIONS ACCT BYPASS=1 METHOD=GEAR
.END
