BICMOS INVERTER PULLDOWN CIRCUIT

VSS 2 0 0V

VIN 3 2 0V (PULSE 0.0V 4.2V 0NS 1NS 1NS 9NS 20NS)

M1  8 3 5 11 M_NMOS_1 W=4U L=1U
VD  4 8 0V
VBK 11 2 0V

Q1  10 7 9   M_NPNS AREA=8
VC  4 10 0V
VB  5 7 0V
VE  9 2 0V

CL  4 6 1PF
VL  6 2 0V

.IC V(10)=5.0V V(7)=0.0V 
.TRAN 0.1NS 5NS 0NS 0.1NS
.PLOT TRAN I(VIN)

.INCLUDE BICMOS.LIB

.OPTIONS ACCT BYPASS=1
.END
