 TIMER 555
 * https://www.electro-tech-online.com/threads/spice-and-555-timer.5806/
 .SUBCKT UA555  32 30 19 23 33 1  21
    *           TR O  R  F  TH D  V
    *
    * Taken from the Fairchild data book (1982) page 9-3
    *SYM=UA555
    *DWG=C:\SPICE\555\UA555.DWG
    Q4 25 2 3 QP
    Q5 0 6 3 QP
    Q6 6 6 8 QP
    R1 9 21 4.7K
    R2 3 21 830
    R3 8 21 4.7K
    Q7 2 33 5 QN
    Q8 2 5 17 QN
    Q9 6 4 17 QN
    Q10 6 23 4 QN
    Q11 12 20 10 QP
    R4 10 21 1K
    Q12 22 11 12 QP
    Q13 14 13 12 QP
    Q14 0 32 11 QP
    Q15 14 18 13 QP
    R5 14 0 100K
    R6 22 0 100K
    R7 17 0 10K
    Q16 1 15 0 QN
    Q17 15 19 31 QP
    R8 18 23 5K
    R9 18 0 5K
    R10 21 23 5K
    Q18 27 20 21 QP
    Q19 20 20 21 QP
    R11 20 31 5K
    D1 31 24 DA
    Q20 24 25 0 QN
    Q21 25 22 0 QN
    Q22 27 24 0 QN
    R12 25 27 4.7K
    R13 21 29 6.8K
    Q23 21 29 28 QN
    Q24 29 27 16 QN
    Q25 30 26 0 QN
    Q26 21 28 30 QN
    D2 30 29 DA
    R14 16 15 100
    R15 16 26 220
    R16 16 0 4.7K
    R17 28 30 3.9K
    Q3 2 2 9 QP
    .MODEL DA D (RS=40 IS=1.0E-14 CJO=1PF)
    .MODEL QP PNP (BF=20 BR=0.02 RC=4 RB=25 IS=1.0E-14 VA=50 NE=2)
    + CJE=12.4P VJE=1.1 MJE=.5 CJC=4.02P VJC=.3 MJC=.3 TF=229P TR=159N)
    .MODEL QN NPN (IS=5.07F NF=1 BF=100 VAF=161 IKF=30M ISE=3.9P NE=2
    + BR=4 NR=1 VAR=16 IKR=45M RE=1.03 RB=4.12 RC=.412 XTB=1.5
    + CJE=12.4P VJE=1.1 MJE=.5 CJC=4.02P VJC=.3 MJC=.3 TF=229P TR=959P)
 .ENDS

    **********
    * Sample Test Circuit for the LM555 Timer: Astable Mode
    * The LM555 timer model is designed for low frequency
    * applications, up to 100Hz.
    .INCLUDE TLC555.LIB
    .TRAN 10u 100MS
    .OPTIONS RELTOL=.0001
    .SAVE  v(16) v(13) v(17)
    .SAVE  v(1) v(4) v(3)

    V2 2 0 5
    VReset res 0 DC 0 PULSE(0 5 1u 1u 1u 30m 50m)

    R3 2 3 1k
    R4 3 4 5k
    C3 4 0 0.5u ; 0.15u
    X2 4  1  res  6  4  3  2 ua555
*      TR O  R    F  TH D  V
    RA 2 17 1k ; 5k
    RB 17 16 5k ; 3k
    C 16 0 0.5u ; 0.15u
    RL 2 13 1k
    X1 16    15   16   res   13  17   2   0   TLC555
*      THRES CONT TRIG RESET OUT DISC VCC GND

    .control
    if $?batchmode
    else
      run
      plot v(16) v(13) v(17) v(1)+6 v(4)+6 v(3)+6
    end
    .endc

    .END
