** PMOSFET: Benchmarking Implementation of BSIM4.3.0 by Jane Xi 05/09/2003.

** Circuit Description **
m1 2 1 0 0 p1 L=0.09u W=10.0u rgeoMod=1
*+SA=0.5u SB=20u geomod=0 sd=0.1u
vgs 1 0 -1.2
vds 2 0 -1.2

.dc vds 0 -1.2 -0.02 vgs -0.3 -1.2 -0.3

.options Temp=100.0
.print dc v(1) i(vds)

.include modelcard.pmos 
.end
