* Param-example
.param amplitude= 1V

.subckt myfilter in out rval=100k  cval=100nF
Ra in p1   {2*rval}
Rb p1 out  {2*rval}
C1 p1 0    {2*cval}
Ca in p2   {cval}
Cb p2 out  {cval}
R1 p2 0    {rval}
.ends myfilter

X1 input output myfilter rval=1k cval=1n
V1 input 0 AC {amplitude}

.end
