psp nch output
*
vd  d 0 dc 0.1
vg  g 0 dc 0.0
vs  s 0 dc 0.0
vb  b 0 dc 0.0
m1  d g s b nch
+l=1.0e-06
+w=10.0e-06
+sa=0.0e+00
+sb=0.0e+00
+absource=1.0e-12
+lssource=1.0e-06
+lgsource=1.0e-06
+abdrain=1.0e-12
+lsdrain=1.0e-06
+lgdrain=1.0e-06
+mult=1.0e+00
*
.option temp=21
.control
dc vd 0 3.5 0.05 vg 0.5 3 0.5
plot abs(i(vd))
plot abs(i(vb)) ylog ylimit 1e-12 1e-03
.endc
*
.model nch nmos level=45
+type=1.0e+00
+tr=21.0e+00
+swigate=0.0e+00
+swimpact=1.0e+00
+swgidl=0.0e+00
+swjuncap=0.0e+00
+lvaro=0.0e+00
+lvarl=0.0e+00
+lvarw=0.0e+00
+lap=0.0e+00
+wvaro=0.0e+00
+wvarl=0.0e+00
+wvarw=0.0e+00
+wot=0.0e+00
+vfbo=-1.0e+00
+vfbl=0.0e+00
+vfbw=0.0e+00
+vfblw=0.0e+00
+stvfbo=500.0e-06
+stvfbl=0.0e+00
+stvfbw=0.0e+00
+stvfblw=0.0e+00
+toxo=2.0e-09
+nsubo=300.0e+21
+nsubw=0.0e+00
+wseg=10.0e-09
+npck=1.0e+24
+npckw=0.0e+00
+wsegp=10.0e-09
+lpck=10.0e-09
+lpckw=0.0e+00
+vnsubo=0.0e+00
+nslpo=50.0e-03
+dnsubo=0.0e+00
+npo=100.0e+24
+npl=0.0e+00
+qmc=1.0e+00
+cto=0.0e+00
+ctl=0.0e+00
+ctlexp=1.0e+00
+ctw=0.0e+00
+toxovo=2.0e-09
+lov=0.0e+00
+novo=50.0e+24
+fol1=0.0e+00
+fol2=0.0e+00
+cfl=0.0e+00
+cflexp=2.0e+00
+cfw=0.0e+00
+cfbo=0.0e+00
+uo=50.0e-03
+fbet1=0.0e+00
+fbet1w=0.0e+00
+lp1=10.0e-09
+lp1w=0.0e+00
+fbet2=0.0e+00
+lp2=10.0e-09
+betw1=0.0e+00
+betw2=0.0e+00
+wbet=1.0e-09
+stbeto=1.0e+00
+stbetl=0.0e+00
+stbetw=0.0e+00
+stbetlw=0.0e+00
+mueo=500.0e-03
+muew=0.0e+00
+stmueo=0.0e+00
+themuo=1.5e+00
+stthemuo=1.5e+00
+cso=0.0e+00
+csw=0.0e+00
+stcso=0.0e+00
+xcoro=0.0e+00
+xcorl=0.0e+00
+xcorw=0.0e+00
+xcorlw=0.0e+00
+stxcoro=0.0e+00
+rsw1=2.5e+03
+rsw2=0.0e+00
+strso=1.0e+00
+rsbo=0.0e+00
+rsgo=0.0e+00
+thesato=0.0e+00
+thesatl=50.0e-03
+thesatlexp=1.0e+00
+thesatw=0.0e+00
+stthesato=1.0e+00
+stthesatl=0.0e+00
+stthesatw=0.0e+00
+stthesatlw=0.0e+00
+thesatbo=0.0e+00
+thesatgo=0.0e+00
+axo=18.0e+00
+axl=400.0e-03
+alpl=500.0e-06
+alplexp=1.0e+00
+alpw=0.0e+00
+alp1l1=0.0e+00
+alp1lexp=500.0e-03
+alp1l2=0.0e+00
+alp1w=0.0e+00
+alp2l1=0.0e+00
+alp2lexp=0.5e+00
+alp2l2=0.0e+00
+alp2w=0.0e+00
+vpo=50.0e-03
+a1o=1.0e+00
+a1l=0.0e+00
+a1w=0.0e+00
+a2o=10.0e+00
+sta2o=0.0e+00
+a3o=1.0e+00
+a3l=0.0e+00
+a3w=0.0e+00
+a4o=0.0e+00
+a4w=0.0e+00
+gcoo=0.0e+00
+iginvlw=0.0e+00
+igovw=0.0e+00
+stigo=2.0e+00
+gc2o=375.0e-03
+gc3o=63.0e-03
+chibo=3.1e+00
+agidlw=0.0e+00
+bgidlo=41.0e+00
+stbgidlo=0.0e+00
+cgidlo=0.0e+00
+cgbovl=0.0e+00
+cfrw=0.0e+00
+nfalw=80.0e+21
+nfblw=30.0e+06
+nfclw=0.0e+00
+saref=1.0e-06
+sbref=1.0e-06
+wlod=0.0e+00
+kuo=0.0e+00
+kvsat=0.0e+00
+tkuo=0.0e+00
+lkuo=0.0e+00
+wkuo=0.0e+00
+pkuo=0.0e+00
+llodkuo=0.0e+00
+wlodkuo=0.0e+00
+kvtho=0.0e+00
+lkvtho=0.0e+00
+wkvtho=0.0e+00
+pkvtho=0.0e+00
+llodvth=0.0e+00
+wlodvth=0.0e+00
+stetao=0.0e+00
+lodetao=1.0e+00
+trj=21.0e+00
+imax=1.0e+03
+cjorbot=1.0e-03
+cjorsti=1.0e-09
+cjorgat=1.0e-09
+vbirbot=1.0e+00
+vbirsti=1.0e+00
+vbirgat=1.0e+00
+pbot=500.0e-03
+psti=500.0e-03
+pgat=500.0e-03
+phigbot=1.16e+00
+phigsti=1.16e+00
+phiggat=1.16e+00
+idsatrbot=1.0e-12
+idsatrsti=1.0e-18
+idsatrgat=1.0e-18
+csrhbot=100.0e+00
+csrhsti=100.0e-06
+csrhgat=100.0e-06
+xjunsti=100.0e-09
+xjungat=100.0e-09
+ctatbot=100.0e+00
+ctatsti=100.0e-06
+ctatgat=100.0e-06
+mefftatbot=250.0e-03
+mefftatsti=250.0e-03
+mefftatgat=250.0e-03
+cbbtbot=1.0e-12
+cbbtsti=1.0e-18
+cbbtgat=1.0e-18
+fbbtrbot=1.0e+09
+fbbtrsti=1.0e+09
+fbbtrgat=1.0e+09
+stfbbtbot=-1.0e-03
+stfbbtsti=-1.0e-03
+stfbbtgat=-1.0e-03
+vbrbot=10.0e+00
+vbrsti=10.0e+00
+vbrgat=10.0e+00
+pbrbot=4.0e+00
+pbrsti=4.0e+00
+pbrgat=4.0e+00
+dta=0.0e+00

.end
