BICMOS 3-STAGE AMPLIFIER
*** IN GRAY & MEYER, 3RD ED. P.266, PROB. 3.12, 8.19

VDD 1 0 5.0V
VSS 2 0 0.0V

*** VOLTAGE INPUT
*VIN 13 0 0.0V AC 1V
*CIN 13 3 1UF

*** CURRENT INPUT
IIN 3 0 0.0 AC 1.0

M1  4 3 2 2 M_NMOS_1 W=300U L=1U
M2  7 7 2 2 M_NMOS_1 W=20U  L=1U

Q1  6 5 4   M_NPNS AREA=40
Q2  5 5 7   M_NPNS AREA=40
Q3  1 6 8   M_NPNS AREA=40

RL1 1 4     1K
RL2 1 6     10K
RB1 1 5     10K
RL3 8 2     1K
RF1 3 8     30K

*** NUMERICAL MODEL LIBRARY ***
.INCLUDE BICMOS.LIB

.AC DEC 10 100KHZ 100GHZ
.PLOT AC VDB(8)

.OPTIONS ACCT BYPASS=1 KEEPOPINFO
.END
