MOS 1 output

m1 d g s b n1 W=40u L=0.8u
.model n1 nmos vt0=1.2

vd d 0 1
vg g 0 1
vs s 0 0
vb b 0 0

.dc vd 0 5 0.1 vg 0 5 1

.control
run
plot vs#branch
.endc

.end
