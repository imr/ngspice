BICMOS INVERTER PULLUP CIRCUIT

VDD 1 0 5.0V
VSS 2 0 0.0V

VIN 3 0 0.75V

VC  1 11 0.0V
VB  5 15 0.0V

Q1  11 15 4 M_NPNS   AREA=8
M1  5 3 1 1 M_PMOS_1 W=10U L=1U

CL  4 0 5.0PF

.IC V(4)=0.75V V(5)=0.0V

.INCLUDE BICMOS.LIB

.TRAN 0.5NS 4.0NS
.PRINT TRAN V(3) V(4)

.OPTION ACCT BYPASS=1
.END
