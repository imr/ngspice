* Random noise test
* internal noise source

* one over f
VNOI1 1 0 DC 0 TRNOISE(0n 1n 1.7 1n)
VNOI2 2 0 DC 0 TRNOISE(0n 1n 1.4 1n)
VNOI3 3 0 DC 0 TRNOISE(0n 1n 1.0 1n)
VNOI4 4 0 DC 0 TRNOISE(0n 1n 0.5 1n)
* white
VNOI5 5 0 DC 0 TRNOISE(1n 1n 0 0)
* both
VNOI6 6 0 DC 0 TRNOISE(1n 1n 1 1n)

* 250000 sample points
.tran 1n 250u

.control
run
plot v(1) v(2) v(3) v(4) v(5) v(6)
plot v(1) v(2) v(3) v(4) v(5) v(6) xlimit 102.0u 102.01u ylimit -3n 3n
linearize
fft v(1) v(2) v(3) v(4) v(5) v(6)
plot mag(v(1)) mag(v(2)) mag(v(3)) mag(v(4)) mag(v(5)) loglog xlimit 1e3 1e9
plot mag(v(6)) loglog xlimit 1e3 1e9
.endc

.end
 
