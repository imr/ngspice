ex3a, check lib processing

I1    7 0  -1mA
X1    7 0  sub1_in_lib

Vcheck1  7 check1  1.0V

I2    9 0  -1mA
X2    9 0  sub2_in_lib

Vcheck2  9 check2  2.0V

.lib 'ex3.lib' MOS

.control
op

let n_pass = 0

echo "Note: v(check1) = $&v(check1)"
echo "Note: v(check2) = $&v(check2)"

if abs(v(check1)) <= 1e-9
    let n_pass = n_pass + 1
else
    echo "ERROR: Test 1 failed"
end


if abs(v(check2)) <= 1e-9
    let n_pass = n_pass + 1
else
    echo "ERROR: Test 2 failed"
end


if n_pass = 2
    echo "INFO: ok"
    quit 0
end

echo ERROR: $&n_pass of 2 tests passed
quit 1

.endc

.end
