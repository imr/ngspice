4 STAGE RTL INVERTER CHAIN

VIN 1 0 DC 0V PWL 0NS 0V 1NS 5V
VCC 12 0 DC 5.0V
RC1 12 3 2.5K
RB1 1 2 8K
Q1 3 2 0 QMOD AREA = 100P
RB2 3 4 8K
RC2 12 5 2.5K
Q2 5 4 0 QMOD AREA = 100P
RB3 5 6 8K
RC3 12 7 2.5K
Q3 7 6 0 QMOD AREA = 100P
RB4 7 8 8K
RC4 12 9 2.5K
Q4 9 8 0 QMOD AREA = 100P

.PRINT TRAN V(3) V(5) V(9)
.TRAN 1E-9 10E-9

.MODEL QMOD NBJT LEVEL=1
+ X.MESH NODE=1  LOC=0.0
+ X.MESH NODE=61 LOC=3.0
+ REGION NUM=1 MATERIAL=1
+ MATERIAL NUM=1 SILICON NBGNN=1E17 NBGNP=1E17
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+ DOPING UNIF N.TYPE CONC=1E17 X.L=0.0 X.H=1.0
+ DOPING UNIF P.TYPE CONC=1E16 X.L=0.0 X.H=1.5
+ DOPING UNIF N.TYPE CONC=1E15 X.L=0.0 X.H=3.0
+ MODELS BGNW SRH CONCTAU AUGER CONCMOB FIELDMOB
+ OPTIONS BASE.LENGTH=1.0 BASE.DEPTH=1.25

.OPTION ACCT BYPASS=1
.END
