DIODE BRIDGE RECTIFIER

VLINE 3 4 0.0V SIN 0V 10V 60HZ
VGRND 2 0 0.0V 
D1 3 1 M_PN AREA=100
D2 4 1 M_PN AREA=100
D3 2 3 M_PN AREA=100
D4 2 4 M_PN AREA=100
RL 1 2 1.0K

.MODEL M_PN NUMD LEVEL=1
+ ***************************************
+ *** ONE-DIMENSIONAL NUMERICAL DIODE ***
+ ***************************************
+ OPTIONS DEFA=1P
+ X.MESH LOC=0.0 N=1
+ X.MESH LOC=30.0 N=201
+ DOMAIN   NUM=1 MATERIAL=1
+ MATERIAL NUM=1 SILICON
+ MOBILITY MAT=1 CONCMOD=CT FIELDMOD=CT
+ DOPING GAUSS P.TYPE CONC=1E20 X.L=0.0  X.H=0.0 CHAR.L=1.0
+ DOPING UNIF  N.TYPE CONC=1E14 X.L=0.0  X.H=30.0
+ DOPING GAUSS N.TYPE CONC=5E19 X.L=30.0  X.H=30.0 CHAR.L=2.0 
+ MODELS BGN ^AVAL SRH AUGER CONCTAU CONCMOB FIELDMOB
+ METHOD AC=DIRECT

.OPTION ACCT BYPASS=1 METHOD=GEAR
.TRAN 0.5MS 50MS
.PRINT TRAN I(VLINE)
.END
