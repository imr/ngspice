** Operational Amplifier (AC): Benchmarking Implementation of BSIM4.7.0 by Mohan V. Dunga 12/13/2006.

M1 bias1 1 cm cm N1 L=0.09u W=10u
M2 bias2 in2 cm cm N1 L=0.09u W=10u
M3 vdd bias1 bias1 vdd P1 L=0.09u W=2u
M4 bias2 bias1 vdd vdd P1 L=0.09u W=2u

m5 cm bias vss vss N1 L=0.09u W=2u
mbias bias bias vss vss N1 L=0.09u W=2u
rbias 0 bias 195k

m6 8 bias vss vss N1 L=0.09u W=2u
m7 8 bias2 vdd out N1 L=0.09u W=2u

Cfb bias2 8 2p

Vid 1 c 0 ac 0.1
eid in2 c 1 c -1
vic c 0 dc 0
vss vss 0 -1.8
Vdd vdd 0 1.8 

.option noacct
.ac dec 10 100 100Meg 
.print ac vdb(8)

.include modelcard.nmos
.include modelcard.pmos

.end
