scope-1, subckt scopes
* (exec-spice "ngspice -b %s" t)

* ----

i1001_t  n1001_t 0  -1mA
x1001_t  n1001_t 0  sub1

v1001_g  n1001_g 0  2.0V

* ----

i1002_t  n1002_t 0  -1mA
x1002_t  n1002_t 0  sub2

v1002_g  n1002_g 0  1.0V

* ----

.subckt  sub1  n1 n2
.subckt  sub   n1 n2
R1   n1 n2   4k
.ends
X1   n1 n2  sub
R1   n1 n2  4k
.ends

.subckt  sub2  n1 n2
.subckt  sub   n1 n2
R1   n1 n2   2k
.ends
X1   n1 n2  sub
R1   n1 n2  2k
.ends


.control

define mismatch(a,b,err) abs(a-b)>err

op

let total_count = 0
let fail_count = 0

let tests = 1001 + vector(2)

foreach n $&tests
  set n_test = "n{$n}_t"
  set n_gold = "n{$n}_g"
  if mismatch(v($n_test), v($n_gold), 1e-9)
    let v_test = v($n_test)
    let v_gold = v($n_gold)
    echo "ERROR, test failure, v($n_test) = $&v_test but should be $&v_gold"
    let fail_count = fail_count + 1
  end
  let total_count = total_count + 1
end

if fail_count > 0
  echo "ERROR: $&fail_count of $&total_count tests failed"
  quit 1
else
  echo "INFO: $&fail_count of $&total_count tests failed"
  quit 0
end

.endc

.end
