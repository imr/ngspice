CMOS RING OSCILLATOR - 1UM DEVICES

VDD 1 0 5.0V
VSS 2 0 0.0V

X1 1 2 3 4 INV
X2 1 2 4 5 INV
X3 1 2 5 6 INV
X4 1 2 6 7 INV
X5 1 2 7 8 INV
X6 1 2 8 9 INV
X7 1 2 9 3 INV

.IC V(3)=0.0V V(4)=2.5V V(5)=5.0V
+   V(6)=0.0V V(7)=5.0V V(8)=0.0V V(9)=5.0V

.SUBCKT INV 1   2   3   4
*           VDD VSS VIN VOUT
M1  14 13 15 16 M_PMOS_1 W=6.0U
M2  24 23 25 26 M_NMOS_1 W=3.0U

VGP 3 13 0.0V
VDP 4 14 0.0V
VSP 1 15 0.0V
VBP 1 16 0.0V

VGN 3 23 0.0V
VDN 4 24 0.0V
VSN 2 25 0.0V
VBN 2 26 0.0V
.ENDS INV

.INCLUDE BICMOS.LIB

.TRAN 0.1NS 1NS
.PRINT TRAN V(3) V(4) V(5)

.OPTIONS ACCT BYPASS=1 METHOD=GEAR
.END
