VOLTAGE CONTROLLED OSCILLATOR

RC1 7 5 1K
RC2 7 6 1K

Q5 7 7 5 QMOD AREA = 100P
Q6 7 7 6 QMOD AREA = 100P

Q3 7 5 2 QMOD AREA = 100P
Q4 7 6 1 QMOD AREA = 100P

IB1 2 0 .5MA
IB2 1 0 .5MA
CB1 2 0 1PF
CB2 1 0 1PF

Q1 5 1 3 QMOD AREA = 100P
Q2 6 2 4 QMOD AREA = 100P

C1 3 4 .1UF 

IS1 3 0 DC 2.5MA PULSE 2.5MA 0.5MA 0 1US 1US 50MS
IS2 4 0 1MA
VCC 7 0 10

.MODEL QMOD NBJT LEVEL=1
+ X.MESH NODE=1  LOC=0.0
+ X.MESH NODE=61 LOC=3.0
+ REGION NUM=1 MATERIAL=1
+ MATERIAL NUM=1 SILICON NBGNN=1E17 NBGNP=1E17
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+ DOPING UNIF N.TYPE CONC=1E17 X.L=0.0 X.H=1.0
+ DOPING UNIF P.TYPE CONC=1E16 X.L=0.0 X.H=1.5
+ DOPING UNIF N.TYPE CONC=1E15 X.L=0.0 X.H=3.0
+ MODELS BGNW SRH CONCTAU AUGER CONCMOB FIELDMOB
+ OPTIONS BASE.LENGTH=1.0 BASE.DEPTH=1.25

.OPTION ACCT BYPASS=1 
.TRAN 3US 600US 0 3US
.PRINT TRAN V(4)
.END
