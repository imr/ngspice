* A fairy tale process deck
* Good for education and examples
* Not good for silicon!
* PTM 90nm NMOS
 
.model  nch  nmos  level = 54

+version = 4.5          binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 1          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0          

+tnom    = 27           toxe    = '2.05e-9-(6E-11*(agauss(0,1,3)))'      toxp    = '1.4e-9-(6E-11*(agauss(0,1,3)))'       toxm    = 2.05e-9   
+epsrox  = 3.9          wint    = 5e-009       lint    = 7.5e-009   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 2.05e-9   
+xl      = '-40e-9-(1E-9*(agauss(0,1,3)))'
+vth0    = '0.397-(0.025*(agauss(0,1,3)))'
+k1      = 0.4          k2      = 0.01         k3      = 0          
+k3b     = 0            w0      = 2.5e-006     dvt0    = 1            dvt1    = 2       
+dvt2    = -0.032       dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 0.1          minv    = 0.05         voffl   = 0            dvtp0   = 1.2e-009     
+dvtp1   = 0.1          lpe0    = 0            lpeb    = 0            xj      = 2.8e-008   
+ngate   = 2e+020       ndep    = 1.94e+018    nsd     = 2e+020       phin    = 0          
+cdsc    = 0.0002       cdscb   = 0            cdscd   = 0            cit     = 0          
+voff    = -0.13        nfactor = 1.7          eta0    = 0.0074       etab    = 0          
+vfb     = -0.55        u0      = 0.0547       ua      = 6e-010       ub      = 1.2e-018     
+uc      = -3e-011      vsat    = 113760       a0      = 1.0          ags     = 1e-020     
+a1      = 0            a2      = 1            b0      = -1e-020      b1      = 0          
+keta    = 0.04         dwg     = 0            dwb     = 0            pclm    = 0.06       
+pdiblc1 = 0.001        pdiblc2 = 0.001        pdiblcb = -0.005       drout   = 0.5        
+pvag    = 1e-020       delta   = 0.01         pscbe1  = 8.14e+008    pscbe2  = 1e-007     
+fprout  = 0.2          pdits   = 0.08         pditsd  = 0.23         pditsl  = 2.3e+006   
+rsh     = 5            rdsw    = 180          rsw     = 90           rdw     = 90        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 0          
+prwb    = 6.8e-011     wr      = 1            alpha0  = 0.074        alpha1  = 0.005      
+beta0   = 30           agidl   = 0.0002       bgidl   = 2.1e+009     cgidl   = 0.0002     
+egidl   = 0.8          

+aigbacc = 0.012        bigbacc = 0.0028       cigbacc = 0.002     
+nigbacc = 1            aigbinv = 0.014        bigbinv = 0.004        cigbinv = 0.004      
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.012        bigc    = 0.0028     
+cigc    = 0.002        aigsd   = 0.012        bigsd   = 0.0028       cigsd   = 0.002     
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1          

+xrcrg1  = 12           xrcrg2  = 5          
+cgso    = 1.9e-010     cgdo    = 1.9e-010     cgbo    = 2.56e-011    cgdl    = 2.653e-10     
+cgsl    = 2.653e-10    ckappas = 0.03         ckappad = 0.03         acde    = 1          
+moin    = 15           noff    = 0.9          voffcv  = 0.02       

+kt1     = -0.11        kt1l    = 0            kt2     = 0.022        ute     = -1.5       
+ua1     = 4.31e-009    ub1     = 7.61e-018    uc1     = -5.6e-011    prt     = 0          
+at      = 33000      

+fnoimod = 1            tnoimod = 0          

+jss     = 0.0001       jsws    = 1e-011       jswgs   = 1e-010       njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 1            cjs     = 0.0005       mjs     = 0.5          pbsws   = 1          
+cjsws   = 5e-010       mjsws   = 0.33         pbswgs  = 1            cjswgs  = 3e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.005        tcj     = 0.001      
+tpbsw   = 0.005        tcjsw   = 0.001        tpbswg  = 0.005        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          

+dmcg    = 0e-006       dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0.0e-008     xgw     = 0e-007       xgl     = 0e-008     

+rshg    = 0.4          gbmin   = 1e-010       rbpb    = 5            rbpd    = 15         
+rbps    = 15           rbdb    = 15           rbsb    = 15           ngcon   = 1          

* PTM 90nm PMOS
 
.model  pch  pmos  level = 54

+version = 4.5          binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 1          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0          

+tnom    = 27           toxe    = '2.15e-009-(6E-11*(agauss(0,1,3)))'    toxp    = '1.4e-009-(6E-11*(agauss(0,1,3)))'     toxm    = 2.15e-009   
+epsrox  = 3.9          wint    = 5e-009       lint    = 7.5e-009   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 2.15e-009   
+xl      = '-40e-9-(1E-9*(agauss(0,1,3)))'
+vth0    = '-0.339-(0.025*(agauss(0,1,3)))'
+k1      = 0.4          k2      = -0.01        k3      = 0          
+k3b     = 0            w0      = 2.5e-006     dvt0    = 1            dvt1    = 2       
+dvt2    = -0.032       dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 0.1          minv    = 0.05         voffl   = 0            dvtp0   = 1e-009     
+dvtp1   = 0.05         lpe0    = 0            lpeb    = 0            xj      = 2.8e-008   
+ngate   = 2e+020       ndep    = 1.43e+018    nsd     = 2e+020       phin    = 0          
+cdsc    = 0.000258     cdscb   = 0            cdscd   = 6.1e-008     cit     = 0          
+voff    = -0.126       nfactor = 1.7          eta0    = 0.0074       etab    = 0          
+vfb     = 0.55         u0      = 0.00711      ua      = 2.0e-009     ub      = 0.5e-018     
+uc      = -3e-011      vsat    = 70000        a0      = 1.0          ags     = 1e-020     
+a1      = 0            a2      = 1            b0      = 0            b1      = 0          
+keta    = -0.047       dwg     = 0            dwb     = 0            pclm    = 0.12       
+pdiblc1 = 0.001        pdiblc2 = 0.001        pdiblcb = 3.4e-008     drout   = 0.56       
+pvag    = 1e-020       delta   = 0.01         pscbe1  = 8.14e+008    pscbe2  = 9.58e-007  
+fprout  = 0.2          pdits   = 0.08         pditsd  = 0.23         pditsl  = 2.3e+006   
+rsh     = 5            rdsw    = 200          rsw     = 100          rdw     = 100        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 3.22e-008  
+prwb    = 6.8e-011     wr      = 1            alpha0  = 0.074        alpha1  = 0.005      
+beta0   = 30           agidl   = 0.0002       bgidl   = 2.1e+009     cgidl   = 0.0002     
+egidl   = 0.8          

+aigbacc = 0.012        bigbacc = 0.0028       cigbacc = 0.002     
+nigbacc = 1            aigbinv = 0.014        bigbinv = 0.004        cigbinv = 0.004      
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.69         bigc    = 0.0012     
+cigc    = 0.0008       aigsd   = 0.0087       bigsd   = 0.0012       cigsd   = 0.0008     
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1 
         
+xrcrg1  = 12           xrcrg2  = 5          
+cgso    = 1.8e-010     cgdo    = 1.8e-010     cgbo    = 2.56e-011    cgdl    = 2.653e-10
+cgsl    = 2.653e-10    ckappas = 0.03         ckappad = 0.03         acde    = 1
+moin    = 15           noff    = 0.9          voffcv  = 0.02

+kt1     = -0.11        kt1l    = 0            kt2     = 0.022        ute     = -1.5       
+ua1     = 4.31e-009    ub1     = 7.61e-018    uc1     = -5.6e-011    prt     = 0          
+at      = 33000      

+fnoimod = 1            tnoimod = 0          

+jss     = 0.0001       jsws    = 1e-011       jswgs   = 1e-010       njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 1            cjs     = 0.0005       mjs     = 0.5          pbsws   = 1          
+cjsws   = 5e-010       mjsws   = 0.33         pbswgs  = 1            cjswgs  = 3e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.005        tcj     = 0.001      
+tpbsw   = 0.005        tcjsw   = 0.001        tpbswg  = 0.005        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          

+dmcg    = 0e-006       dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0.0e-008     xgw     = 0e-007       xgl     = 0e-008     

+rshg    = 0.4          gbmin   = 1e-010       rbpb    = 5            rbpd    = 15         
+rbps    = 15           rbdb    = 15           rbsb    = 15           ngcon   = 1          

*****3.3V IO MOS******

.model  nio  nmos  level = 54

+version = 4.0          binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 1          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0


+tnom    = 27           
+toxe    = '7e-9-(2E-10*(agauss(0,1,3)))'      
+toxp    = '7e-9-(2E-10*(agauss(0,1,3)))'       toxm    = 7e-9   
+epsrox  = 3.9           wint    = 4.5e-008       lint    = 2e-008   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 7e-9   
+xl      = '-2e-8-(2E-8*(agauss(0,1,3)))'
+vth0    = '-0.55-(0.015*(agauss(0,1,3)))'



+k1      = 0.7          k2      = -0.03        k3      = 0          
+k3b     = 0            w0      = 0            dvt0    = 0            dvt1    = 2       
+dvt2    = -0.032       dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 0.5          minv    = 0.05         voffl   = 0            dvtp0   = 0     
+dvtp1   = 0.1          lpe0    = 0            lpeb    = 0            xj      = 2.8e-008   
+ngate   = 4.5e+021     ndep    = 1.74e+017    nsd     = 1e+020       phin    = 0.1          
+cdsc    = 0.0002       cdscb   = 0            cdscd   = 0            cit     = 0          
+voff    = -0.1         nfactor = 1            eta0    = 0.05         etab    = -0.16          
+vfb     = -0.55        u0      = 0.02         ua      = 8e-010       ub      = 7.8e-019     
+uc      = -2e-011      vsat    = 7600         a0      = 1.4          ags     = 0.21     
+a1      = 0            a2      = 1            b0      = -1e-020      b1      = 0          
+keta    = -0.014       dwg     = 0            dwb     = 0            pclm    = 0.36       
+pdiblc1 = 0            pdiblc2 = 0.00014      pdiblcb = 0            drout   = 0.5        
+pvag    = 1e-020       delta   = 0.006        pscbe1  = 8.14e+008    pscbe2  = 2e-005     
+fprout  = 0.2          pdits   = 0.08         pditsd  = 0.23         pditsl  = 2.3e+006   
+rsh     = 10           rdsw    = 540          rsw     = 270          rdw     = 270        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 1          
+prwb    = 6.8e-011     wr      = 1            alpha0  = 0.001        alpha1  = 1      
+beta0   = 40           agidl   = 2e-10        bgidl   = 1.7e+009     cgidl   = 0.7     
+egidl   = 0.48                   


+aigbacc = 0.4          bigbacc = 0.054        cigbacc = 0.075     
+nigbacc = 1            aigbinv = 0.35         bigbinv = 0.03         cigbinv = 0.006      
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.4          bigc    = 0.06     
+cigc    = 0.075        aigsd   = 0.4          bigsd   = 0.05         cigsd   = 0.075     
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1


+xrcrg1  = 12           xrcrg2  = 1          
+cgso    = 7.3e-011     cgdo    = 7.3e-011     cgbo    = 0            cgdl    = 2e-10     
+cgsl    = 2e-10        ckappas = 0.03         ckappad = 0.03         acde    = 0.5          
+moin    = 5            noff    = 1.63         voffcv  = -0.02       

+kt1     = -0.345       kt1l    = 0            kt2     = -0.035       ute     = -0.35       
+ua1     = 3.6e-10      ub1     = -1.6e-018    uc1     = -3e-011      prt     = 0          
+at      = 170000      

+fnoimod = 1            tnoimod = 0 


+jss     = 1.5e-007     jsws    = 5.3e-014     jswgs   = 4.3e-014     njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 0.75         cjs     = 0.00122      mjs     = 0.33         pbsws   = 1          
+cjsws   = 1.56e-011    mjsws   = -0.11        pbswgs  = 0.75         cjswgs  = 2.7e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.0017       tcj     = 0.0009      
+tpbsw   = 0.0002       tcjsw   = 0.0003       tpbswg  = 0.001        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          

+dmcg    = 1.0e-007     dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0.0e-008     xgw     = 0e-007       xgl     = 0e-008     

+rshg    = 0.1          gbmin   = 1e-012       rbpb    = 50           rbpd    = 50         
+rbps    = 50           rbdb    = 50           rbsb    = 50           ngcon   = 1




.model  pio  pmos  level = 54

+version = 4.0          binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 1          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0


+tnom    = 27           
+toxe    = '7e-9-(2E-10*(agauss(0,1,3)))'      
+toxp    = '7e-9-(2E-10*(agauss(0,1,3)))'      toxm    = 7e-9   
+epsrox  = 3.9           wint    = 9.5e-008     lint    = 6e-008   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 7e-9   
+xl      = '-2e-8-(2E-8*(agauss(0,1,3)))'
+vth0    = '-0.65-(0.015*(agauss(0,1,3)))'



+k1      = 0.7          k2      = -0.03        k3      = 0          
+k3b     = 0            w0      = 0            dvt0    = 0            dvt1    = 2       
+dvt2    = -0.032       dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 0.5          minv    = 0.05         voffl   = 0            dvtp0   = 0     
+dvtp1   = 0.1          lpe0    = 0            lpeb    = 0            xj      = 2.8e-008   
+ngate   = 4.5e+021     ndep    = 1.74e+017    nsd     = 1e+020       phin    = 0.1          
+cdsc    = 0.0002       cdscb   = 0            cdscd   = 0            cit     = 0          
+voff    = -0.1         nfactor = 1            eta0    = 0.05         etab    = -0.16          
+vfb     = -0.55        u0      = 0.011        ua      = 8e-010       ub      = 7.8e-019     
+uc      = -2e-011      vsat    = 7600         a0      = 1.4          ags     = 0.21     
+a1      = 0            a2      = 1            b0      = -1e-020      b1      = 0          
+keta    = -0.014       dwg     = 0            dwb     = 0            pclm    = 0.36       
+pdiblc1 = 0            pdiblc2 = 0.00014      pdiblcb = 0            drout   = 0.5        
+pvag    = 1e-020       delta   = 0.006        pscbe1  = 8.14e+008    pscbe2  = 2e-005     
+fprout  = 0.2          pdits   = 0.08         pditsd  = 0.23         pditsl  = 2.3e+006   
+rsh     = 10           rdsw    = 540          rsw     = 270          rdw     = 270        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 1          
+prwb    = 6.8e-011     wr      = 1            alpha0  = 0.001        alpha1  = 1      
+beta0   = 40           agidl   = 2e-10        bgidl   = 1.7e+009     cgidl   = 0.7     
+egidl   = 0.48                   


+aigbacc = 0.4          bigbacc = 0.054        cigbacc = 0.075     
+nigbacc = 1            aigbinv = 0.35         bigbinv = 0.03         cigbinv = 0.006      
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.4          bigc    = 0.06     
+cigc    = 0.075        aigsd   = 0.4          bigsd   = 0.05         cigsd   = 0.075     
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1


+xrcrg1  = 12           xrcrg2  = 1          
+cgso    = 7.3e-011     cgdo    = 7.3e-011     cgbo    = 0            cgdl    = 2e-10     
+cgsl    = 2e-10        ckappas = 0.03         ckappad = 0.03         acde    = 0.5          
+moin    = 5            noff    = 1.63         voffcv  = -0.02       

+kt1     = -0.345       kt1l    = 0            kt2     = -0.035       ute     = -0.35       
+ua1     = 3.6e-10      ub1     = -1.6e-018    uc1     = -3e-011      prt     = 0          
+at      = 170000      

+fnoimod = 1            tnoimod = 0 






*****resistors******
.model hrp r
+TC1R     = -6E-04     	    TC2R     = 1.08E-06        
+DW       = '6E-08'         DLR  = -6.5E-07
+TNOM     = 27              RSH      = '1000-(200*(agauss(0,1,3)))'

.model lrp r
*poly resistor
+TC1R     = 2.69E-03      TC2R     = -2.65E-06
+DW = '2.5E-08-(1.01E-08*(agauss(0,1,3)))'
+TNOM     = 27            RSH      = '10-(2.2*(agauss(0,1,3)))'


.model mrp r 
*poly resistor  
+TC1R     = 1.2E-04      TC2R     = -9E-08
+DW       = '4E-08-(8E-09*(agauss(0,1,3)))'       DLR = -1.5E-07 
+TNOM     = 27            RSH      = '100-(17.689*(agauss(0,1,3)))'

*****BJT*****
.model pnp PNP
+LEVEL    = 1                   
+VAF      = 700                 IKF      = 7.2E-03          
+ISE      = 7E-17               NE       = 1.5                BR       = 4E-03          
+NR       = 1                   VAR      = 80                 IKR      = 4E-03           
+ISC      = 1.5E-16             NC       = 1.5                RB       = 55             
+IRB      = 1.6E-03             RBM      = 5.1346             RE       = 1.0                 
+RC       = 10.0                XTI      = 3.0                EG       = 1.16                
+TREF     = 27                  NKF      = 0.5                TLEV     = 0
+TLEVC    = 1                   XTB      = 0.00               TBF1     = 4E-03          
+TBF2     = 3.9E-06             TBR1     = -2.3E-03           TBR2     = 1.6E-05            
+TIKF1    = -2.4E-03            TIKF2    = -1.12E-05          TNF1     = 1.1E-06           
+TNF2     = -5.74E-07           TNR1     = 2.5E-05            TNR2     = -1.3E-06         
+TRB1     = 1.6E-03             TRB2     = 7E-06            
+TNE1     = -10E-04             TNE2     = -1.2E-05         
+TRM1     = 0                   TRM2     = 0                         
+CTC      = 2E-03               CTE      = 9E-04              
+VJE      = 0.8                 MJE      = 0.3                 SUBS     = 1
+VJC      = 0.6                 MJC      = 0.45                                  
+TVJC     = 1.8E-03             TVJE     = 1.7E-03
+IS       = '6.4E-18+(1.28E-18*(agauss(0,1,3)))'  
+BF       = '0.9+(1.2E-01*(agauss(0,1,3)))'             
+NF       = '1.02-(0.008*(agauss(0,1,3)))'
+CJC      = '9E-14-(4.59E-15*(agauss(0,1,3)))'
+CJE      = '1E-13-(6.13E-15*(agauss(0,1,3)))'
