.title KiCad schematic
.include "./models/TLV9002.LIB"
Vsignal1 Vin GND dc 2.5 ac 1
Vcc1 Vcc GND 5
R1 Vin Net-_R1-Pad2_ 1000
R2 Vout Net-_R1-Pad2_ 1meg
R3 Vcc Net-_R3-Pad2_ 10k
R4 Net-_R3-Pad2_ GND 10k
XU1 Net-_R3-Pad2_ Net-_R1-Pad2_ Vcc GND Vout TLV9002
.save @vsignal1[i]
.save @vcc1[i]
.save @r1[i]
.save @r2[i]
.save @r3[i]
.save @r4[i]
.save V(Net-_R1-Pad2_)
.save V(Net-_R3-Pad2_)
.save V(Vcc)
.save V(Vin)
.save V(Vout)
.ac dec 10 100m 20k

*.options NOOPITER GMINSTEPS=0
*.options  RELTOL=1e-3 VNTOL=1u PIVTOL=1e-11

.control
optran 0 0 0 100n 10u 0
run
plot db(Vout)
set units=degrees
plot ph(Vout)
.endc

.end
