*not per Fra

.include ./models/16nm_HP.pm

*.model p1_ra relmodel level=1 h_cut=b nts=c m_star=f w=g tau_0=h beta=i tau_e=j beta1=k
*.model p1_ra relmodel level=1 tau_0=5e-12 beta=0.746
.model p1_ra relmodel level=1 type=1
.appendmodel p1_ra pmos

.meas tran delay_LH trig v(in) val=0.5 fall=1 targ v(out) val=0.5 rise=1
.meas tran delay_HL trig v(in) val=0.5 rise=1 targ v(out) val=0.5 fall=1

Mp1 OUT IN Vdd Vdd pmos L=22n W=44n
Mn1 OUT IN 0 0     nmos L=22n W=22n

Cl out 0 10f

Valim Vdd 0 0.7
*Vin IN 0 pwl(0 0 10n 0 11n 1 60n 1 61n 0 110n 0 111n 1 160n 1 161n 0 210n 0 211n 1 260n 1
*+            261n 0 310n 0 311n 1 360n 1 361n 0 410n 0 411n 1 460n 1 461n 0 510n 0 511n 1 560n 1
*+            561n 0 610n 0 611n 1 660n 1 661n 0 710n 0 711n 1 760n 1 761n 0 810n 0 811n 1 860n 1
*+            861n 0)
*Vin IN 0 pwl(0 0 0.5n 0 0.501n 1 1n 1 1.01n 0 1.5n 0 1.501n 1 2n 1 2.01n 0 2.5n 0 2.501n 1 3n 1 3.01n 0 3.5n 0 3.501n 1 4n 1
*+            4.01n 0 4.5n 0 4.501n 1 5n 1 5.01n 0 5.5n 0 5.501n 1 6n 1 6.01n 0 6.5n 0 6.501n 1 7n 1 7.01n 0 7.5n 0 7.501n 1 8n 1
*+            8.01n 0 8.5n 0 8.501n 1 9n 1 9.01n 0 9.5n 0 9.501n 1 10n 1)
Vin IN 0 pwl(0 0 2n 0 2.01n 0.7 4n 0.7 4.01n 0 6n 0 6.01n 0.7 8n 0.7 8.01n 0 10n 0 10.01n 0.7 12n 0.7 12.01n 0 14n 0 14.01n 0.7 16n 0.7
+            16.01n 0 18n 0 18.01n 0.7 20n 0.7 20.01n 0 22n 0 22.01n 0.7 24n 0.7 24.01n 0 26n 0 26.01n 0.7 28n 0.7 28.01n 0 30n 0 30.01n 0.7 32n 0.7
+            32.01n 0 34n 0 34.01n 0.7 36n 0.7 36.01n 0 38n 0 38.01n 0.7 40n 0.7 40.01n 0 42n 0 42.01n 0.7 44n 0.7 44.01n 0 46n 0 46.01n 0.7 48n 0.7)
*Vin IN 0 pwl(0 0 10n 0)
*Vin IN 0 pwl(0 1 10n 1)

.relan 315360000 10p 48n
.tran 10p 48n

.control 
  run
.endc
