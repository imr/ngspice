* Mesa Test
* Taken from macspice3f4

z1 3 2 0 mesmod l=1u w=150u
vgs 2 0 dc 0
vds 1 0 dc 0
vids 1 3 dc 0

.model mesmod nmf level=3 rdi=2.7 rsi=2.7 mu=0.2 m=2.2 vto=-2.04
+ eta=1.5 lambda=0.04 tc=0.001 sigma0=0.02 vsigma=0.1 vsigmat=1.37
+ delta=5 beta=0.0085

.options noacct

.dc vds 0 4 0.05 vgs -1.5 0.5 0.5
.print vids#branch

.end

