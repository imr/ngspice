* MESA1 transient test 
* Taken from macspice3f4
* 
* This netlist shows convergence problems in ngspice

rd 1 3 10k
z1 3 2 0 mesa1 l=1u w=20u
vgs 2 0 dc 0 pulse(-3 0 0 0.5n 0.5n 2n 4n)
vdd  1 0 5v
.model mesa1 nmf(level=2 rd=31 rs=31)

.options noacct
.dc vgs -2 0 0.02
.tran 0.1n 5n
.print tran v(2) v(3)

.print 
