vdmos model test

mn1 d s g b IRFZ48Z

.model IRFZ48Z VDMOS ( Rg = 1.77 Vto=4 Rd=1.85m Rs=0.0m Rb=3.75m Kp=25 Cgdmax=2.1n Cgdmin=0.05n Cgs=1.8n Cjo=0.55n Is=2.5p tt=20n mfg=International_Rectifier Vds=55 Ron=8.6m Qg=43n)

mn2 d2 s2 g2 b2 SUM110P04-05
.MODEL SUM110P04-05 VDMOS(KP=80 RS=0.002 RD=0.001 RG=3.0 VTO=-3.3 LAMBDA=0.05 CGDMAX=7n CGDMIN=800p CGS=9n TT=100n a=0.55 IS=1.5E-08 N=1.35 RB=0.001 m=0.774 Vj=1.59 Cjo=3nF PCHAN)

.end