  ADDER - 4 BIT ALL-74HC00-GATE BINARY ADDER WITH AUTOMATIC BRIDGING
  * behavioral gate description
  * Automatic A/D insertion using bi-directional bridges

* Override the default bridges and force use of the bidi_bridges with
* directions controlled by inputs.

.control
pre_set auto_bridge_d_out =
+ ( ".model auto_bridge_out bidi_bridge(out_high=%g)"
+   "auto_bridge_out%d [ %s ] [ %s ] [ force_out ] auto_bridge_out"  1 )
pre_set auto_bridge_d_in =
+ ( ".model auto_bridge_in bidi_bridge(in_low='%g/2' in_high='%g/2')"
+   "auto_bridge_in%d [ %s ] [ %s ] [ force_in ] auto_bridge_in" 1  )
.endc

*** SUBCIRCUIT DEFINITIONS
.include 74HCng_auto.lib
.param vcc=3 tripdt=6n

aup force_in pullup
.model pullup d_pullup
adown force_out pulldown
.model pulldown d_pulldown

.include ../adder_common.inc

.END
