rca3040 ckt - rca 3040 wideband amplifier
.options noacct
.ac dec 10 1 10ghz
.dc vin -0.25 0.25 0.005
.tran 2.0ns 200ns
vin 1 0 sin(0 0.1 50meg 0.5ns) ac 1
vcc     2       0       15.0
vee     3       0       -15.0
rs1     30      1       1k
rs2     31      0       1k
r1      5       3       4.8k
r2      6       3       4.8k
r3      9       3       811
r4      8       3       2.17k
r5      8       0       820
r6      2       14      1.32k
r7      2       12      4.5k
r8      2       15      1.32k
r9      16      0       5.25k
r10     17      0       5.25k
q1      2       30      5       qnl
q2      2       31      6       qnl
q3      10      5       7       qnl
q4      11      6       7       qnl
q5      14      12      10      qnl
q6      15      12      11      qnl
q7      12      12      13      qnl
q8      13      13      0       qnl
q9      7       8       9       qnl
q10     2       15      16      qnl
q11     2       14      17      qnl
.model qnl npn level=1 bf=80 rb=100 ccs=2pf tf=0.3ns tr=6ns cje=3pf
+ cjc=2pf va=50
.end
