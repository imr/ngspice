VDMOS output

m1 d g s s IXTP6N100D2
m2 d g s2 s2 IXTP6N100D2_2

*.model dmod d  is=10n rs=0.05

* LTSPICE model parameters
*.MODEL IXTP6N100D2 VDMOS(KP=2.9 RS=0.1 RD=1.3 RG=1 VTO=-2.7 LAMBDA=0.03 CGDMAX=3000p CGDMIN=2p CGS=2915p TT=1371n a=1 IS=2.13E-08 N=1.564 RB=0.0038 m=0.548 *Vj=0.1 Cjo=3200pF subthres=2.5m)

* equivalent ngspice model parameters
.MODEL IXTP6N100D2 VDMOS(KP=2.9 RS=0.1 RD=1.3 RG=1 VTO=-2.7 LAMBDA=0.03 CGDMAX=3000p CGDMIN=2p CGS=2915p TT=1371n a=1 IS=2.13E-08 N=1.564 RB=0.0038 m=0.548 Vj=0.1 Cjo=3200pF subslope=43m subshift=-25m)

vd d 0 -0.6
vg g 0 -2.3
vs s 0 0

.control
dc  vg -3.1 -2.1 0.01 vd 0.2 1 0.2
plot vs#branch
plot vs#branch ylog
dc  vd 0 5 0.01 vg -3.2 -2 0.2
plot vs#branch
.endc

.end
