ECL INVERTER
*** (FROM MEINERZHAGEN ET AL.)

VCC 1 0 0.0V
VEE 2 0 -5.2V

VIN 3 0 -1.25V
VRF 4 0 -1.25V

*** INPUT STAGE
Q1 5 3 9 M_NPNS AREA=8
Q2 6 4 9 M_NPNS AREA=8
R1 1 5 662
R2 1 6 662
R3 9 2 2.65K

*** OUTPUT BUFFERS
Q3 1 5 7 M_NPNS AREA=8
Q4 1 6 8 M_NPNS AREA=8
R4 7 2 4.06K
R5 8 2 4.06K

*** MODEL LIBRARY
.INCLUDE BICMOS.LIB

.DC VIN -2.00 0.001 0.05
.PLOT DC V(7) V(8)

.OPTIONS ACCT BYPASS=1
.END
