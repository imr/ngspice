BICMOS INVERTER PULLUP CIRCUIT

VDD 1 0 5.0V
VSS 2 0 0.0V

VIN 3 0 0.75V

VC  1 11 0.0V
VB  5 15 0.0V

Q1  11 15 4 M_NPN  AREA=4
M1  5 3 1 1 M_PMOS W=20U L=2U AD=30P AS=30P PD=21U PS=21U

CL  4 0 5.0PF

.IC V(4)=0.75V V(5)=0.0V

.MODEL M_PMOS PMOS VTO=-0.8 UO=250 TOX=25N NSUB=5E16
+ UCRIT=10K UEXP=.15 VMAX=50K NEFF=2 XJ=.02U
+ LD=.15U CGSO=.1N CGDO=.1N CJ=.12M MJ=0.5
+ CJSW=0.3N MJSW=0.5 LEVEL=2

.MODEL M_NPN NBJT LEVEL=2
+ TITLE TWO-DIMENSIONAL NUMERICAL POLYSILICON EMITTER BIPOLAR TRANSISTOR
+ $ SINCE ONLY HALF THE DEVICE IS SIMULATED, DOUBLE THE UNIT WIDTH TO GET
+ $ 1.0 UM EMITTER.
+ OPTIONS DEFW=2.0U
+ OUTPUT STATISTICS
+ 
+ X.MESH W=2.0 H.E=0.02 H.M=0.5 R=2.0
+ X.MESH W=0.5 H.S=0.02 H.M=0.2 R=2.0
+ 
+ Y.MESH L=-0.2 N=1
+ Y.MESH L= 0.0 N=5
+ Y.MESH W=0.10 H.E=0.004 H.M=0.05  R=2.5
+ Y.MESH W=0.15 H.S=0.004 H.M=0.02  R=2.5
+ Y.MESH W=1.05 H.S=0.02  H.M=0.1   R=2.5
+
+ DOMAIN NUM=1 MATERIAL=1 X.L=2.0 Y.H=0.0
+ DOMAIN NUM=2 MATERIAL=2 X.H=2.0 Y.H=0.0
+ DOMAIN NUM=3 MATERIAL=3 Y.L=0.0
+ MATERIAL NUM=1 POLYSILICON
+ MATERIAL NUM=2 OXIDE
+ MATERIAL NUM=3 SILICON
+
+ ELEC NUM=1 X.L=0.0  X.H=0.0  Y.L=1.1  Y.H=1.3
+ ELEC NUM=2 X.L=0.0  X.H=0.5  Y.L=0.0  Y.H=0.0
+ ELEC NUM=3 X.L=2.0  X.H=3.0  Y.L=-0.2 Y.H=-0.2
+
+ DOPING GAUSS N.TYPE CONC=3E20 X.L=2.0 X.H=3.0 Y.L=-0.2 Y.H=0.0
+ + CHAR.L=0.047 LAT.ROTATE
+ DOPING GAUSS P.TYPE CONC=5E18 X.L=0.0 X.H=5.0 Y.L=-0.2 Y.H=0.0
+ + CHAR.L=0.100 LAT.ROTATE
+ DOPING GAUSS P.TYPE CONC=1E20 X.L=0.0 X.H=0.5 Y.L=-0.2 Y.H=0.0
+ + CHAR.L=0.100 LAT.ROTATE RATIO=0.7
+ DOPING UNIF  N.TYPE CONC=1E16 X.L=0.0 X.H=5.0 Y.L=0.0 Y.H=1.3
+ DOPING GAUSS N.TYPE CONC=5E19 X.L=0.0 X.H=5.0 Y.L=1.3 Y.H=1.3
+ + CHAR.L=0.100 LAT.ROTATE
+
+ METHOD AC=DIRECT ITLIM=10
+ MODELS BGN SRH AUGER CONCTAU CONCMOB FIELDMOB

.TRAN 0.5NS 4.0NS
.PRINT TRAN V(3) V(4)

.OPTION ACCT BYPASS=1
.END
