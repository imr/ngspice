OpAmp Test

vddp vp 0 3
vddn vn 0 -3

*vin in 0 0

* OPA171 IN+ IN- VCC VEE OUT
.include OPA171.txt

Xopmap 0 ino vp vn outo OPA171

*Xopmap 0 ino outo vp vn CLC409
Rin in ino 1k
Rfb ino outo 3k

*.dc vin -1 1 0.1

vin in 0 DC 0 PULSE(-0.5 0.5 2uS 200NS 200NS 5uS 10uS)
.tran 100n 10u

.control
run
plot v(in) v(outo)
.endc


*
*   This is a Very Wide band, Low Distortion Monolithic
*   Current Feedback Op Amp.
*
* Version 1, Rev. A, Date 04-09-92, By RRS
*
* Connections: Non-Inverting Input
*              | Inverting Input
*              | | Output
*              | | | +Vcc
*              | | | | -Vcc
*              | | | | |
.SUBCKT CLC409 3 2 6 7 4
*
* DC BIAS MIRROR
*
R1 7 4 28K
R2 7 9 271
R3 10 4 335
*
G1 7 11 POLY(2) 7 9 7 4 0 3.15M 21.5U
C3 11 0 128F
*
G2 14 4 POLY(1) 10 4 0 2.95M
C4 14 0 104F
*
* INPUT VOLTAGE BUFFER
*
E1 3 17 POLY(1) 35 0 1.0M 1.673
C6 17 0 1.00P
*
Q1 10 17 12 QINP
D3 11 12 DY
Q2 9 17 13 QINN
D4 13 14 DY
*
G3 2 0 POLY(1) 36 0 0 9.282M
C10 2 0 2.9P
*
D5 22 2 DY
Q3 21 11 22 QINN
D6 2 23 DY
Q4 24 14 23 QINP
*
* CURRENT MIRROR GAIN BLOCKS
*
R10 7 20 640
V1 20 21 1.9
C8 21 28 294F
G4 7 28 POLY(1) 7 20 0 4.3M
R15 7 28 102K
C13 28 0 641F
D1 28 26 DX
V3 7 26 1.65
G6 7 30 POLY(1) 7 20 0 2.74M
C15 30 0 676F
*
R13 25 4 640
V2 24 25 1.85
C12 24 29 294F
G5 29 4 POLY(1) 25 4 0 4.5M
R16 29 4 761K
C14 29 0 312F
D2 27 29 DX
V4 27 4 1.55
G7 31 4 POLY(1) 25 4 0 6.74M
C16 31 0 330F
*
* OUTPUT STAGE AND COMPENSATION CAPACITORS
*
R14 28 29 45.0
Q5 4 29 30 QOUTP1
Q6 7 28 31 QOUTN1
*
C9 21 33 .935P
C11 24 33 .935P
C17 33 0 4.00P
R19 33 6 10
*
Q7 7 30 33 QOUTN2
Q8 4 31 33 QOUTP2
*
* NOISE BLOCKS
*
R20 35 0 122
R21 35 0 122
*
R22 36 0 122
R23 36 0 122
*
* MODELS
*
.MODEL DX D TT=200N
.MODEL DY D IS=0.166F
*
.MODEL QINN NPN
+ IS =0.166f    BF =3.239E+02 NF =1.000E+00 VAF=8.457E+01
+ IKF=2.462E-02 ISE=2.956E-17 NE =1.197E+00 BR =3.719E+01
+ NR =1.000E+00 VAR=1.696E+00 IKR=3.964E-02 ISC=1.835E-19
+ NC =1.700E+00 RB =118       IRB=0.000E+00 RBM=65.1
+ RC =2.645E+01 CJE=1.632E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.948E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=5.955E-02 PTF=0.000E+00 CJC=1.720E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=589m     TR =4.212E-10 CJS=629f
+ MJS=0         KF =2.000E-12 AF =1.000E+00 FC =9.765E-01
*
.MODEL QOUTN1 NPN
+ IS =3.954E-16 BF =3.239E+02  NF =1.000E+00 VAF=8.457E+01
+ IKF=4.590E-02 ISE=5.512E-17  NE =1.197E+00 BR =3.719E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=7.392E-02 ISC=3.087E-19
+ NC =1.700E+00 RB =3.645E+01  IRB=0.000E+00 RBM=8.077E+00
+ RE =3.010E-01 RC =2.702E+01  CJE=2.962E-13
+ MJE=4.950E-01 TF =1.904E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=1.110E-01 PTF=0.000E+00  CJC=2.846E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.562E-01 TR =5.832E-10 CJS=5.015E-13
+ VJS=5.723E-01 MJS=4.105E-01  KF =2.000E-12 AF =1.000E+00
+ FC =9.765E-01
*
.MODEL QOUTN2 NPN
+ IS =9.386E-16 BF =3.239E+02 NF =1.000E+00 VAF=8.457E+01
+ IKF=1.089E-01 ISE=1.308E-16 NE =1.197E+00 BR =3.956E+01
+ NR =1.000E+00 VAR=1.696E+00 IKR=7.392E-02 ISC=1.378E-18
+ NC =1.700E+00 RB =65.4      IRB=0.000E+00 RBM=1.683E+00
+ RC =1.857E+01 CJE=7.030E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.875E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=2.635E-01 PTF=0.000E+00 CJC=6.172E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=860m     TR =1.069E-09 CJS=1.028E-12
+ VJS=5.723E-01 MJS=4.105E-01 KF =2.000E-12 AF =1.000E+00
+ FC =9.765E-01
*
.MODEL QINP PNP
+ IS =0.166f    BF =7.165E+01 NF =1.000E+00 VAF=2.000E+01
+ IKF=1.882E-02 ISE=6.380E-16 NE =1.366E+00 BR =1.833E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=1.321E-01 ISC=3.666E-18
+ NC =1.634E+00 RB =78.8      IRB=0.000E+00 RBM=57.6
+ RC =3.739E+01 CJE=1.588E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.156E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=5.084E-02 PTF=0.000E+00 CJC=2.725E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=741m     TR =7.500E-11 CJS=515f
+ MJS=0         KF =2.000E-12 AF =1.000E+00 FC =8.803E-01
*
.MODEL QOUTP1 PNP
+ IS =2.399E-16 BF =7.165E+01  NF =1.000E+00 VAF=3.439E+01
+ IKF=3.509E-02 ISE=1.190E-15  NE =1.366E+00 BR =1.900E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=2.464E-01 ISC=6.745E-18
+ NC =1.634E+00 RB =1.542E+01  IRB=0.000E+00 RBM=4.059E+00
+ RC =4.174E+01 CJE=2.962E-13  VJE=7.975E-01
+ MJE=5.000E-01 TF =3.107E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=9.481E-02 PTF=0.000E+00  CJC=4.508E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.562E-01 TR =9.500E-11 CJS=1.045E-12
+ VJS=6.691E-01 MJS=3.950E-01  KF =2.000E-12 AF =1.000E+00
+ FC =8.803E-01
*
.MODEL QOUTP2 PNP
+ IS =5.693E-16 BF =7.165E+01 NF =1.000E+00 VAF=3.439E+01
+ IKF=8.328E-02 ISE=5.742E-15 NE =1.366E+00 BR =1.923E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=5.848E-01 ISC=1.586E-17
+ NC =1.634E+00 RB =56.5      IRB=0.000E+00 RBM=51.7
+ RC =1.767E+00 CJE=7.030E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.073E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=2.250E-01 PTF=0.000E+00 CJC=9.776E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=923m     TR =1.450E-10 CJS=1.637E-12
+ VJS=6.691E-01 MJS=3.950E-01 KF =2.000E-12 AF =1.000E+00
+ FC =8.803E-01
*
.ENDS CLC409

.end

