A Simple AC Run

.OPTIONS LIST NODE POST TRANS
.OP
.AC DEC 10 1k 1Meg
.PRINT AC V(2)

V1 1 0 DC 0 AC 1 SIN 0 1 1K 0 0 DISTOF1 0 DISTOF2 0
R1 1 2 10k
R2 2 0 10k
C1 2 0 1n

.END
