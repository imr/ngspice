RTL inverter

vin 1 0 dc 1 pwl 0 4 1ns 0
vcc 12 0 dc 5.0
rc1 12 3 2.5k
rb1 1 2 8k
q1 3 2 0 qmod area = 100p

.option acct bypass=1
.tran 0.5n 5n
.print tran v(2) v(3)

.model qmod nbjt level=1
+ x.mesh node=1  loc=0.0
+ x.mesh node=61 loc=3.0
+ region num=1 material=1
+ material num=1 silicon nbgnn=1e17 nbgnp=1e17
+ mobility material=1 concmod=sg fieldmod=sg
+ mobility material=1 elec major
+ mobility material=1 elec minor
+ mobility material=1 hole major
+ mobility material=1 hole minor
+ doping unif n.type conc=1e17 x.l=0.0 x.h=1.0
+ doping unif p.type conc=1e16 x.l=0.0 x.h=1.5
+ doping unif n.type conc=1e15 x.l=0.0 x.h=3.0
+ models bgnw srh conctau auger concmob fieldmob
+ options base.length=1.0 base.depth=1.25

.end
