PUSH-PULL EMITTER FOLLOWER - ONE-DIMENSIONAL MODELS

VCC 1 0  5.0V
VEE 2 0 -5.0V

VIN 3 0  0.0V (SIN 0.0V 0.1V 1KHZ) AC 1
VBU 13 3 0.7V
VBL 3 23 0.7V

RL  4 44  50
VLD 44 0 0V

Q1  5  13 4 M_NPN1D AREA=40
Q2  4  5  1 M_PNP1D AREA=200

Q3  6  23 4 M_PNP1D AREA=100
Q4  4  6  2 M_NPN1D AREA=80

.INCLUDE BICMOS.LIB

.TRAN 0.01MS 1.00001MS 0US 0.01MS
.PLOT TRAN V(4)

.OPTIONS ACCT BYPASS=1 TEMP=26.85OC RELTOL=1E-5
.END
