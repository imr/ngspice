** One-Shot Trigger (Tran): Benchmarking Implementation of BSIM4.0.0 by Weidong Liu 5/16/2000.

Md1 4 in Vdd Vdd  P1 W=3.6u L=1.2u
Md2 4 in 0 0 N1 W=1.8u L=1.2u
c4 4 0 30f
Md3 A 4 Vdd Vdd  P1 W=3.6u L=1.2u
Md4 A 4 0 0 N1 W=1.8u L=1.2u
ca a 0 30f

M1 Anot A Vdd Vdd  P1 W=3.6u L=1.2u
M2 Anot A 0 0 N1 W=1.8u L=1.2u

M3 Bnot in Vdd Vdd  P1 W=3.6u L=1.2u
M4 Bnot in 0 0 N1 W=1.8u L=1.2u

M5 AorBnot 0 Vdd Vdd P1 W=1.8u L=3.6u
M6 AorBnot in 1 0 N1 W=1.8u L=1.2u
M7 1 Anot 0 0 N1 W=1.8u L=1.2u

M8 Lnot 0 Vdd Vdd P1 W=1.8u L=3.6u
M9 Lnot Bnot 2 0 N1 W=1.8u L=1.2u
M10 2 A 0 0 N1 W=1.8u L=1.2u

M11 out 0 Vdd Vdd P1 W=3.6u L=3.6u
M12 out AorBnot 3 0 N1 W=1.8u L=1.2u
M13 3 Lnot 0 0 N1 W=1.8u L=1.2u

Vcc vdd 0 1.8
vin in 0 pulse 0 1.8 1ns .1ns .1ns .8ns 5ns

.include modelcard.nmos
.include modelcard.pmos

.tran 1ns 10ns
.print tran in out
.option post

.end
