4 Stage RTL Inverter Chain

vin 1 0 dc 0v pwl 0ns 0v 1ns 5v
vcc 12 0 dc 5.0v
rc1 12 3 2.5k
rb1 1 2 8k
q1 3 2 0 qmod area = 100p
rb2 3 4 8k
rc2 12 5 2.5k
q2 5 4 0 qmod area = 100p
rb3 5 6 8k
rc3 12 7 2.5k
q3 7 6 0 qmod area = 100p
rb4 7 8 8k
rc4 12 9 2.5k
q4 9 8 0 qmod area = 100p

.print tran v(3) v(5) v(9)
.tran 1e-9 10e-9

.model qmod nbjt level=1
+ x.mesh node=1  loc=0.0
+ x.mesh node=61 loc=3.0
+ region num=1 material=1
+ material num=1 silicon nbgnn=1e17 nbgnp=1e17
+ mobility material=1 concmod=sg fieldmod=sg
+ mobility material=1 elec major
+ mobility material=1 elec minor
+ mobility material=1 hole major
+ mobility material=1 hole minor
+ doping unif n.type conc=1e17 x.l=0.0 x.h=1.0
+ doping unif p.type conc=1e16 x.l=0.0 x.h=1.5
+ doping unif n.type conc=1e15 x.l=0.0 x.h=3.0
+ models bgnw srh conctau auger concmob fieldmob
+ options base.length=1.0 base.depth=1.25

.option acct bypass=1
.end
