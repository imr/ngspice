CMOS RING OSCILLATOR - 2UM DEVICES

VDD 1 0 5.0V
VSS 2 0 0.0V

X1 1 2 3 4 INV
X2 1 2 4 5 INV
X3 1 2 5 6 INV
X4 1 2 6 7 INV
X5 1 2 7 8 INV
X6 1 2 8 9 INV
X7 1 2 9 3 INV

.IC V(3)=0.0V V(4)=2.5V V(5)=5.0V V(6)=0.0V
+ V(7)=5.0V V(8)=0.0V V(9)=5.0V

.SUBCKT INV 1   2   3   4
*           VDD VSS VIN VOUT
M1  14 13 15 16 M_PMOS W=6.0U
M2  24 23 25 26 M_NMOS W=3.0U

VGP 3 13 0.0V
VDP 4 14 0.0V
VSP 1 15 0.0V
VBP 1 16 0.0V

VGN 3 23 0.0V
VDN 4 24 0.0V
VSN 2 25 0.0V
VBN 2 26 0.0V
.ENDS INV

.MODEL M_NMOS NUMOS
+ X.MESH L=0.0 N=1
+ X.MESH L=0.6 N=4
+ X.MESH L=0.7 N=5
+ X.MESH L=1.0 N=7
+ X.MESH L=1.2 N=11
+ X.MESH L=3.2 N=21
+ X.MESH L=3.4 N=25
+ X.MESH L=3.7 N=27
+ X.MESH L=3.8 N=28
+ X.MESH L=4.4 N=31
+
+ Y.MESH L=-.05 N=1
+ Y.MESH L=0.0  N=5
+ Y.MESH L=.05  N=9
+ Y.MESH L=0.3  N=14
+ Y.MESH L=2.0  N=19
+
+ REGION NUM=1 MATERIAL=1 Y.L=0.0
+ MATERIAL NUM=1 SILICON
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+
+ REGION NUM=2 MATERIAL=2 Y.H=0.0 X.L=0.7 X.H=3.7
+ MATERIAL NUM=2 OXIDE
+
+ ELEC NUM=1 X.L=3.8 X.H=4.4	Y.L=0.0 Y.H=0.0
+ ELEC NUM=2 X.L=0.7 X.H=3.7	IY.L=1  IY.H=1
+ ELEC NUM=3 X.L=0.0 X.H=0.6	Y.L=0.0 Y.H=0.0
+ ELEC NUM=4 X.L=0.0 X.H=4.4	Y.L=2.0 Y.H=2.0
+
+ DOPING UNIF P.TYPE CONC=2.5E16 X.L=0.0 X.H=4.4  Y.L=0.0 Y.H=2.0
+ DOPING UNIF P.TYPE CONC=1E16   X.L=0.0 X.H=4.4  Y.L=0.0 Y.H=0.05
+ DOPING UNIF N.TYPE CONC=1E20   X.L=0.0 X.H=1.1  Y.L=0.0 Y.H=0.2
+ DOPING UNIF N.TYPE CONC=1E20   X.L=3.3 X.H=4.4  Y.L=0.0 Y.H=0.2
+
+ MODELS CONCMOB FIELDMOB BGN SRH CONCTAU
+ METHOD AC=DIRECT ONEC
+ OUTPUT ^ALL.DEBUG

.MODEL M_PMOS NUMOS
+ X.MESH L=0.0 N=1
+ X.MESH L=0.6 N=4
+ X.MESH L=0.7 N=5
+ X.MESH L=1.0 N=7
+ X.MESH L=1.2 N=11
+ X.MESH L=3.2 N=21
+ X.MESH L=3.4 N=25
+ X.MESH L=3.7 N=27
+ X.MESH L=3.8 N=28
+ X.MESH L=4.4 N=31
+
+ Y.MESH L=-.05 N=1
+ Y.MESH L=0.0  N=5
+ Y.MESH L=.05  N=9
+ Y.MESH L=0.3  N=14
+ Y.MESH L=2.0  N=19
+
+ REGION NUM=1 MATERIAL=1 Y.L=0.0
+ MATERIAL NUM=1 SILICON
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+
+ REGION NUM=2 MATERIAL=2 Y.H=0.0 X.L=0.7 X.H=3.7
+ MATERIAL NUM=2 OXIDE
+
+ ELEC NUM=1 X.L=3.8 X.H=4.4	Y.L=0.0 Y.H=0.0
+ ELEC NUM=2 X.L=0.7 X.H=3.7	IY.L=1  IY.H=1
+ ELEC NUM=3 X.L=0.0 X.H=0.6	Y.L=0.0 Y.H=0.0
+ ELEC NUM=4 X.L=0.0 X.H=4.4	Y.L=2.0 Y.H=2.0
+
+ DOPING UNIF N.TYPE CONC=1E16   X.L=0.0 X.H=4.4  Y.L=0.0 Y.H=2.0
+ DOPING UNIF P.TYPE CONC=3E16   X.L=0.0 X.H=4.4  Y.L=0.0 Y.H=0.05
+ DOPING UNIF P.TYPE CONC=1E20   X.L=0.0 X.H=1.1  Y.L=0.0 Y.H=0.2
+ DOPING UNIF P.TYPE CONC=1E20   X.L=3.3 X.H=4.4  Y.L=0.0 Y.H=0.2
+
+ MODELS CONCMOB FIELDMOB BGN SRH CONCTAU
+ METHOD AC=DIRECT ONEC
+ OUTPUT ^ALL.DEBUG

.TRAN 0.1NS 5.0NS
.PRINT V(4)
.OPTIONS ACCT BYPASS=1 METHOD=GEAR
.END
