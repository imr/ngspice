* delta sigma modulator 
* first order, continuous time

.subckt mod1 ainp ainn dclk ddffq ddffqb
* integrator and summer
Ri1 ainn inintn 500
Rf1 adffq inintn 500
Cint1 outintp inintn 1n
.IC v(outintp) = 0 v(inintp) = 0
*
Rshunt1 outintp 0 100Meg
Rshunt2 initn 0 100Meg
*
Ri2 ainp inintp 500
Rf2 adffqb inintp 500
Cint2 outintn inintp 1n
.IC v(outintn) = 0 v(inintn) = 0
*
Rshunt3 outintn 0 100Meg
Rshunt4 inintp 0 100Meg
*
aint %vd(inintp inintn) %vd(outintp outintn) amp
.model amp gain ( in_offset =0.0 gain =100000
+ out_offset = 0)

* latched comparator (code model or B source, analog in, digital out)
*acomp %vd(outintp outintn) acompout limit5
*.model limit5 limit(in_offset=0 gain=100000 out_lower_limit=-1.0
*+ out_upper_limit=1.0 limit_range=0.10 fraction=FALSE)
*
BComp acompout 0 V = (V(outintp) - V(outintn)) >= 0 ? 1 : -1
*
abridge2 [acompout] [dcompout] adc_buff
.model adc_buff adc_bridge(in_low = 0 in_high = 0)
*
* D flip flop: data clk set reset out nout
adff1 dcompout dclk ds drs ddffq ddffqb flop2
.model flop2 d_dff(clk_delay = 1e-9 set_delay = 1.0e-9
+ reset_delay = 1.0e-9 ic = 0 rise_delay = 1.0e-9
+ fall_delay = 1e-9)

abridge1 [ddffq ddffqb dclk] [adffq adffqb aclk] dac1
.model dac1 dac_bridge(out_low = -1 out_high = 1 out_undef = 0
+ input_load = 5.0e-12

.ends mod1
