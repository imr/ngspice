** PMOSFET: Benchmarking Implementation of BSIM4.4.0 by Jane Xi 01/30/2004.

** Circuit Description **
m1 2 1 0 b p1 L=0.09u W=10.0u rgeoMod=1
vgs 1 0 -1.2
vds 2 0 -1.2
vbs b 0 0.0

*.dc vds 0 -1.2 -0.02 vgs 0 -1.2 -0.3
.dc vbs -0.5 2 0.02
*.options Temp=300

.print dc v(1) i(vds)

.include modelcard.pmos 
.end
