prog1-4.cir
 
*** analysis type ***
.tran .01us 10us
v1 1 0 DC 1.0
v2 2 0 DC 0.0

.model d_osc1 d_osc (cntl_array=[-1.0 0.0 1.0 2.0] 
+                    freq_array=[1.0e6 1.0e6 4.0e6 4.0e6]
+                    rise_delay=1.0e-6 fall_delay=2.0e-6)

a1 1 clk1 d_osc1 
a2 2 clk2 d_osc1 

ap0_4 null clk1 null [q1 q2 q3 q4] proc0
.model proc0 d_process (process_file="graycode" process_params=["none"])

ap1_4 [clk2] clk1 null [o1 o2 o3 o4] proc1
.model proc1 d_process (process_file="prog1in4out" process_params=["opt1", "qwerty"])

ap4_1 [o1 o2 o3 o4] clk1 null [zeros] proc2
.model proc2 d_process (process_file="prog4in1out" process_params=["abc", "99"])

ap4_1a [q1 q2 q3 q4] clk1 null [qzeros] proc3
.model proc3 d_process (process_file="prog4in1out")

an1 [o1 ~o2 o3] reseto dand1
.model dand1 d_and(inertial_delay=true rise_delay=1ns fall_delay=50ns)

ap1_4a [clk2] clk1 reseto [b1 b2 b3 b4] proc4
.model proc4 d_process (process_file="prog1in4out")

.control
run
edisplay
eprvcd clk1 clk2  o1 o2 o3 o4 q1 q2 q3 q4 b1 b2 b3 b4 zeros qzeros reseto > prog1-4.vcd
if $oscompiled = 1 | $oscompiled = 8  ; MS Windows
  shell start gtkwave prog1-4.vcd --script nggtk.tcl
else
  shell gtkwave prog1-4.vcd --script nggtk.tcl &
end
quit
.endc
.end






