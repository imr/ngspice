* MLIN test

V1 1 4 PULSE(0 1 1n 10p 10p 980p)
V3 4 0 DC 1
R1 out 2 20.0
V2 2 0 0
R2 in 1 1m
*R3 in ins 1e12
*R4 out outs 1e12
A1 %hd(in 0) %hd(out 0) %vd(in 0) %vd(out 0) MLIN1
.MODEL MLIN1 MLIN(w=1e-3 l=50e-3 er=9.8 h=1e-3 t=35e-6 tand=1e-3 rho=0.022e-6 d=0.15e-6 model=0 disp=0 tranmodel=1)
*A1 %hd(in 0) %hd(out 0) %vd(in 0) %vd(out 0) TLIN1
*.MODEL TLIN1 TLINE(l=100e-3 z=50.0 a=0.0)

.control

*op
*print all

tran 10p 5n

plot v(in) v(out)
plot -i(v1) i(V2)

.endc
