** One-Bit Comparator (Tran): Benchmarking Implementation of BSIM4.7.0 by Mohan V. Dunga 12/13/2006.

M1 Anot A Vdd Vdd  P1 W=3.6u L=0.2u rgeomod=1
M2 Anot A 0 0 N1 W=1.8u L=0.2u rgeomod=1
M3 Bnot B Vdd Vdd  P1 W=3.6u L=0.2u rgeomod=1
M4 Bnot B 0 0 N1 W=1.8u L=0.2u rgeomod=1
M5 AorBnot 0 Vdd Vdd P1 W=1.8u L=3.6u rgeomod=1
M6 AorBnot B 1 0 N1 W=1.8u L=0.2u rgeomod=1
M7 1 Anot 0 0 N1 W=1.8u L=0.2u rgeomod=1
M8 Lnot 0 Vdd Vdd P1 W=1.8u L=3.6u rgeomod=1
M9 Lnot Bnot 2 0 N1 W=1.8u L=0.2u rgeomod=1
M10 2 A 0 0 N1 W=1.8u L=0.2u rgeomod=1
M11 Qnot 0 Vdd Vdd P1 W=3.6u L=3.6u rgeomod=1
M12 Qnot AorBnot 3 0 N1 W=1.8u L=0.2u rgeomod=1
M13 3 Lnot 0 0 N1 W=1.8u L=0.2u rgeomod=1
MQLO 8 Qnot Vdd Vdd  P1 W=3.6u L=0.2u rgeomod=1
MQL1 8 Qnot 0 0 N1 W=1.8u L=0.2u rgeomod=1
MLTO 9 Lnot Vdd Vdd P1 W=3.6u L=0.2u rgeomod=1
MLT1 9 Lnot 0 0 N1 W=1.8u L=0.2u rgeomod=1
CQ Qnot 0 30f
CL Lnot 0 10f

Vdd Vdd 0 1.8
Va A 0  pulse 0 1.8 10ns .1ns .1ns 15ns 30ns
Vb B 0 0

.include modelcard.nmos
.include modelcard.pmos

.tran 1ns 60ns
.option reltol=1e-3 post noacct
.print tran a b v(9) v(8) 

.end
