Component type 283 : 4-bit adder with analog IN/OUT ports

.param vcc=3.2

.subckt 283  a1 a2 a3 a4 b1 b2 b3 b4 c0 sigma1 sigma2 sigma3 sigma4 c4
+     optional: DPWR=$G_DPWR DGND=$G_DGND
+     params: MNTYMXDLY=0 IO_LEVEL=0

U1 BUF $G_DPWR $G_DGND  2 3
+ M1 IOM1 IO_LEVEL=0 MNTYMXDLY=2
U2 AND(2) $G_DPWR $G_DGND  4 5 6
+ M2 IOM2 IO_LEVEL=0 MNTYMXDLY=2
U3 AND(3) $G_DPWR $G_DGND  7 5 8 9
+ M3 IOM3 IO_LEVEL=0 MNTYMXDLY=2
U4 AND(4) $G_DPWR $G_DGND  10 5 8 11 12
+ M4 IOM4 IO_LEVEL=0 MNTYMXDLY=2
U5 AND(5) $G_DPWR $G_DGND  5 8 11 13 14 15
+ M5 IOM5 IO_LEVEL=0 MNTYMXDLY=2
U6 NOR(5) $G_DPWR $G_DGND  3 6 9 12 15 C4
+ M6 IOM6 IO_LEVEL=0 MNTYMXDLY=2
U7 INV $G_DPWR $G_DGND  2 17
+ M7 IOM7 IO_LEVEL=0 MNTYMXDLY=2
U8 AND(2) $G_DPWR $G_DGND  5 17 18
+ M8 IOM8 IO_LEVEL=0 MNTYMXDLY=2
U9 BUF $G_DPWR $G_DGND  4 19
+ M9 IOM9 IO_LEVEL=0 MNTYMXDLY=2
U10 AND(2) $G_DPWR $G_DGND  7 8 20
+ M10 IOM10 IO_LEVEL=0 MNTYMXDLY=2
U11 AND(3) $G_DPWR $G_DGND  10 8 11 21
+ M11 IOM11 IO_LEVEL=0 MNTYMXDLY=2
U12 AND(4) $G_DPWR $G_DGND  8 11 13 14 22
+ M12 IOM12 IO_LEVEL=0 MNTYMXDLY=2
U13 NOR(4) $G_DPWR $G_DGND  19 20 21 22 23
+ M13 IOM13 IO_LEVEL=0 MNTYMXDLY=2
U15 INV $G_DPWR $G_DGND  4 24
+ M15 IOM15 IO_LEVEL=0 MNTYMXDLY=2
U16 AND(2) $G_DPWR $G_DGND  8 24 25
+ M16 IOM16 IO_LEVEL=0 MNTYMXDLY=2
U17 BUF $G_DPWR $G_DGND  7 26
+ M17 IOM17 IO_LEVEL=0 MNTYMXDLY=2
U18 AND(2) $G_DPWR $G_DGND  10 11 27
+ M18 IOM18 IO_LEVEL=0 MNTYMXDLY=2
U19 AND(3) $G_DPWR $G_DGND  11 13 14 28
+ M19 IOM19 IO_LEVEL=0 MNTYMXDLY=2
U21 NOR(3) $G_DPWR $G_DGND  26 27 28 29
+ M21 IOM21 IO_LEVEL=0 MNTYMXDLY=2
U22 INV $G_DPWR $G_DGND  7 30
+ M22 IOM22 IO_LEVEL=0 MNTYMXDLY=2
U23 AND(2) $G_DPWR $G_DGND  11 30 31
+ M23 IOM23 IO_LEVEL=0 MNTYMXDLY=2
U24 BUF $G_DPWR $G_DGND  10 32
+ M24 IOM24 IO_LEVEL=0 MNTYMXDLY=2
U25 AND(2) $G_DPWR $G_DGND  13 14 33
+ M25 IOM25 IO_LEVEL=0 MNTYMXDLY=2
U26 NOR(2) $G_DPWR $G_DGND  32 33 34
+ M26 IOM26 IO_LEVEL=0 MNTYMXDLY=2
U28 INV $G_DPWR $G_DGND  10 35
+ M28 IOM28 IO_LEVEL=0 MNTYMXDLY=2
U29 AND(2) $G_DPWR $G_DGND  13 35 36
+ M29 IOM29 IO_LEVEL=0 MNTYMXDLY=2
U30 INV $G_DPWR $G_DGND  14 37
+ M30 IOM30 IO_LEVEL=0 MNTYMXDLY=2
U32 INV $G_DPWR $G_DGND  C0 14
+ M32 IOM32 IO_LEVEL=0 MNTYMXDLY=2
U33 NAND(2) $G_DPWR $G_DGND  b1 a1 13
+ M33 IOM33 IO_LEVEL=0 MNTYMXDLY=2
U34 NOR(2) $G_DPWR $G_DGND  b1 a1 10
+ M34 IOM34 IO_LEVEL=0 MNTYMXDLY=2
U35 NOR(2) $G_DPWR $G_DGND  B2 A2 7
+ M35 IOM35 IO_LEVEL=0 MNTYMXDLY=2
U36 NAND(2) $G_DPWR $G_DGND  B2 A2 11
+ M36 IOM36 IO_LEVEL=0 MNTYMXDLY=2
U37 NAND(2) $G_DPWR $G_DGND  b3 A3 8
+ M37 IOM37 IO_LEVEL=0 MNTYMXDLY=2
U38 NOR(2) $G_DPWR $G_DGND  b3 A3 4
+ M38 IOM38 IO_LEVEL=0 MNTYMXDLY=2
U39 NOR(2) $G_DPWR $G_DGND  B4 A4 2
+ M39 IOM39 IO_LEVEL=0 MNTYMXDLY=2
U40 NAND(2) $G_DPWR $G_DGND  B4 A4 5
+ M40 IOM40 IO_LEVEL=0 MNTYMXDLY=2
*** U41 STIM(8,44) $G_DPWR $G_DGND  a1 A2 A3 A4 b1 B2 b3 B4
*** + IO_STD IO_LEVEL=0
*** + LABEL=START   0NS INCR BY 11   100NS GOTO START -1 TIMES 
*** U42 STIM(1,1) $G_DPWR $G_DGND  C0
*** + IO_STD IO_LEVEL=0
*** + 0NS 0 
U43 XOR $G_DPWR $G_DGND  18 23 SIGMA4
+ M1 IO_STD IO_LEVEL=0 MNTYMXDLY=2
U44 XOR $G_DPWR $G_DGND  25 29 SIGMA3
+ M1 IO_STD IO_LEVEL=0 MNTYMXDLY=2
U45 XOR $G_DPWR $G_DGND  31 34 SIGMA2
+ M1 IO_STD IO_LEVEL=0 MNTYMXDLY=2
U46 XOR $G_DPWR $G_DGND  36 37 SIGMA1
+ M1 IO_STD IO_LEVEL=0 MNTYMXDLY=2
*
.MODEL M1 UGATE (TPLHTY=3N TPHLTY=2N)
.MODEL IOM1 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M2 UGATE ()
.MODEL IOM2 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M3 UGATE ()
.MODEL IOM3 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M4 UGATE ()
.MODEL IOM4 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M5 UGATE ()
.MODEL IOM5 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M6 UGATE ()
.MODEL IOM6 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M7 UGATE ()
.MODEL IOM7 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M8 UGATE ()
.MODEL IOM8 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M9 UGATE ()
.MODEL IOM9 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M10 UGATE ()
.MODEL IOM10 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M11 UGATE ()
.MODEL IOM11 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M12 UGATE ()
.MODEL IOM12 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M13 UGATE ()
.MODEL IOM13 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M14 UGATE ()
.MODEL IOM14 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M15 UGATE ()
.MODEL IOM15 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M16 UGATE ()
.MODEL IOM16 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M17 UGATE ()
.MODEL IOM17 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M18 UGATE ()
.MODEL IOM18 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M19 UGATE ()
.MODEL IOM19 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M20 UGATE ()
.MODEL IOM20 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M21 UGATE ()
.MODEL IOM21 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M22 UGATE ()
.MODEL IOM22 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M23 UGATE ()
.MODEL IOM23 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M24 UGATE ()
.MODEL IOM24 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M25 UGATE ()
.MODEL IOM25 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M26 UGATE ()
.MODEL IOM26 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M27 UGATE ()
.MODEL IOM27 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M28 UGATE ()
.MODEL IOM28 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M29 UGATE ()
.MODEL IOM29 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M30 UGATE ()
.MODEL IOM30 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M31 UGATE ()
.MODEL IOM31 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M32 UGATE ()
.MODEL IOM32 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M33 UGATE ()
.MODEL IOM33 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M34 UGATE ()
.MODEL IOM34 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M35 UGATE ()
.MODEL IOM35 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M36 UGATE ()
.MODEL IOM36 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M37 UGATE ()
.MODEL IOM37 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M38 UGATE ()
.MODEL IOM38 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M39 UGATE ()
.MODEL IOM39 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
.MODEL M40 UGATE (TPLHTY=4N TPHLTY=6N)
.MODEL IOM40 UIO (INLD=0 OUTLD=0 DRVH=50 DRVL=50 ATOD1="ATOD1" 
+ DTOA1="DTOD1" ATOD2="ATOD2" DTOA2="DTOD2" ATOD3="ATOD3" DTOA3="DTOD3" 
+ ATOD4="ATOD4" DTOA4="DTOD4" TSWLH1=0 TSWLH2=0 TSWLH3=0 TSWLH4=0 
+ TSWHL1=0 TSWHL2=0 TSWHL3=0 TSWHL4=0 DIGPOWER="DIGPOWER")
*** From file C:\MC12\library\DIGIO.LIB
.MODEL IO_STD UIO (
+  DRVH=130 DRVL=130
+  ATOD1="ATOD_STD" ATOD2="ATOD_STD_NX"
+  ATOD3="ATOD_STD" ATOD4="ATOD_STD_NX"
+  DTOA1="DTOA_STD" DTOA2="DTOA_STD"
+  DTOA3="DTOA_STD" DTOA4="DTOA_STD"
+  TSWHL1=3.310NS TSWHL2=3.310NS
+  TSWHL3=3.310NS TSWHL4=3.310NS
+  TSWLH1=2.115NS TSWLH2=2.115NS
+  TSWLH3=2.115NS TSWLH4=2.115NS
+  DIGPOWER="DIGIFPWR")
*
.ends 283

X1 a1 a2 a3 a4 b1 b2 b3 b4 c0 sigma1 sigma2 sigma3 sigma4 c4 283

va1 a1 0 pulse( 0.0 3.2 0ns 0ns 0ns 100ns 200ns )
va2 a2 0 pulse( 3.2 0.0 0ns 0ns 0ns 100ns 200ns )
va3 a3 0 pulse( 0.0 3.2 0ns 0ns 0ns 100ns 200ns )
va4 a4 0 pulse( 3.2 0.0 0ns 0ns 0ns 100ns 200ns )

vb1 b1 0 pulse( 3.2 0.0 0ns 0ns 0ns 100ns 200ns )
vb2 b2 0 pulse( 3.2 0.0 0ns 0ns 0ns 100ns 200ns )
vb3 b3 0 pulse( 3.2 0.0 0ns 0ns 0ns 100ns 200ns )
vb4 b4 0 pulse( 0.0 3.2 0ns 0ns 0ns 100ns 200ns )

vc0 c0 0 pulse( 0.0 3.2 2us )

r1 a1 0 10k
r2 a2 0 10k
r3 a3 0 10k
r4 a4 0 10k
r5 c0 0 10k
r6 c4 0 10k
r10 b1 0 10k
r20 b2 0 10k
r30 b3 0 10k
r40 b4 0 10k
r100 sigma1 0 10k
r200 sigma2 0 10k
r300 sigma3 0 10k
r400 sigma4 0 10k

.tran 1ns 4us
.control
run
listing expand
edisplay
* eprint a4 a3 a2 a1 b4 b3 b2 b1 c0
* eprint sigma4 sigma3 sigma2 sigma1 c4
* save data to input directory
cd $inputdir 
eprvcd a4 a3 a2 a1 b4 b3 b2 b1 c0 sigma4 sigma3 sigma2 sigma1 c4 > ab_ex283.vcd
* plotting the vcd file with GTKWave
if $oscompiled = 1 | $oscompiled = 8  ; MS Windows
  shell start gtkwave ab_ex283.vcd --script nggtk.tcl
else
  if $oscompiled = 7 ; macOS, manual tweaking required (mark, insert, Zoom Fit)
    shell open -a gtkwave ab_ex283.vcd
  else ; Linux and others
    shell gtkwave ab_ex283.vcd --script nggtk.tcl &
  end
end
quit
.endc
.end
