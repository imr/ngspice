Behavioral CMOS 283 : 4-bit adder

*-------------------------------------------------------------74AC283-----
*
* The 74AC283 4-Bit Binary Full Adder with Fast Carry
* (4 Page Fax) Harris Advanced CMOS Logic, File Number 1912
* and Philips Semiconductors High-speed CMOS Logic Data Handbook 
* for the logic diagram, 1994, page 564
* jat 7/26/95

.SUBCKT 74AC283
+ A0 A1 A2 A3 B0 B1 B2 B3 CIN COUT S0 S1 S2 S3
+ OPTIONAL: DPWR=$G_DPWR DGND=$G_DGND
+ PARAMS: MNTYMXDLY=0 IO_LEVEL=0

U1 LOGICEXP(9,5) DPWR DGND
+ A0 A1 A2 A3 B0 B1 B2 B3 CIN 
+ S_0 S_1 S_2 S_3 C_OUT
+ D0_GATE IO_AC
+ MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}
+ LOGIC:
+        S_0 = {A0 ^ B0 ^ CIN}
+        NOR1 = {(A0 | B0) & (CIN | (A0 & B0))}
+        S_1 = {NOR1 ^ A1 ^ B1}
+        NOR2 = {~((~(A1 | B1)) | ((~(A0 | B0)) & (~(A1 & B1))) | 
+          ((~(A1 & B1)) & (~(A0 & B0)) & (~CIN)))}
+        S_2 = {NOR2 ^ A2 ^ B2}
+        AND31 = {(~(A2 & B2)) & (~(A1 & B1)) & (~(A0 & B0)) & (~CIN)}
+        AND32 = {(~(A0 | B0)) & (~(A2 & B2)) & (~(A1 & B1))}
+        AND33 = {(~(A1 | B1)) & (~(A2 & B2))}
+        NOR3 = {~(AND31 | AND32 | AND33 | (~(A2 | B2)))}
+        S_3 = {NOR3 ^ A3 ^ B3}
+        ANDC1 = {(~(A3 & B3)) & (~(A2 & B2)) & (~(A1 & B1)) &
+           (~(A0 & B0)) & (~CIN)}
+        ANDC2 = {(~(A0 | B0)) & (~(A3 & B3)) & (~(A2 & B2)) & (~(A1 & B1))}
+        ANDC3 = {(~(A1 | B1)) & (~(A3 & B3)) & (~(A2 & B2))}
+        ANDC4 = {(~(A2 | B2)) & (~(A3 & B3))}
+        C_OUT = {~(ANDC1 | ANDC2 | ANDC3 | ANDC4 | (~(A3 | B3)))}

U2 PINDLY(5,0,9) DPWR DGND
+ S_0 S_1 S_2 S_3 C_OUT
+ A0 A1 A2 A3 B0 B1 B2 B3 CIN
+ S0 S1 S2 S3 COUT
+ IO_AC
+ MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}
+ BOOLEAN:
+          CARRYIN = {CHANGED(CIN,0)}
+          NUMBER = {CHANGED(A0,0) | CHANGED(A1,0) | CHANGED(A2,0) |
+                    CHANGED(A3,0) | CHANGED(B0,0) | CHANGED(B1,0) |
+                    CHANGED(B2,0) | CHANGED(B3,0)}
+ PINDLY:
+          S0 S1 S2 S3 = {
+             CASE(
+                NUMBER & (TRN_LH | TRN_HL), DELAY(4.7NS,-1,16.5NS),
+                CARRYIN & (TRN_LH | TRN_HL), DELAY(4.5NS,-1,16NS),
+                DELAY(5.7NS,-1,17.5NS))}
+          COUT = {
+             CASE(
+                NUMBER & (TRN_LH | TRN_HL), DELAY(4.5NS,-1,16NS),
+                CARRYIN & (TRN_LH | TRN_HL), DELAY(4.5NS,-1,16NS),
+                DELAY(5.7NS,-1,17.5NS))}

.ENDS 74AC283

X1 a0 a1 a2 a3 b0 b1 b2 b3 cin cout s0 s1 s2 s3 74ac283
a_1 [ a3 a2 a1 a0 b3 b2 b1 b0 cin ] input_vec1
.model input_vec1 d_source(input_file = "ex283.stim")

.tran 0.01ns 2us
.control
run
listing
edisplay
eprint a3 a2 a1 a0 b3 b2 b1 b0 cin
eprint s3 s2 s1 s0 cout
* save data to input directory
cd $inputdir 
eprvcd a3 a2 a1 a0 b3 b2 b1 b0 cin s3 s2 s1 s0 cout > behav-283.vcd
* plotting the vcd file with GTKWave
if $oscompiled = 1 | $oscompiled = 8  ; MS Windows
  shell start gtkwave behav-283.vcd --script nggtk.tcl
else
  shell gtkwave behav-283.vcd --script nggtk.tcl &
end
quit
.endc
.end
