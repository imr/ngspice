*** NDINV * 4
XNDINV1 1 11 12 13 2 100 NDINV
XNDINV2 2 21 22 23 3 100 NDINV
XNDINV3 3 31 32 33 4 100 NDINV
XNDINV4 4 41 42 43 5 100 NDINV

.SUBCKT NDINV 10 11 21 31 41 100
MP11  11 100 100 100   P12L5   L=1.2U W=5U
MP12  11 100 100 100   P12L5   L=1.2U W=5U
MP13  11 100 100 100   P12L5   L=1.2U W=5U
MP14  11  10 100 100   P12L5   L=1.2U W=5U
MN11  11 100  12   0   N10L5   L=1.0U W=5U
MN12  12 100  13   0   N10L5   L=1.0U W=5U
MN13  13 100  14   0   N10L5   L=1.0U W=5U
MN14  14  10   0   0   N10L5   L=1.0U W=5U

MP21  23   0 100 100   P12L5   L=1.2U W=20U
MP22  22  11  23 100   P12L5   L=1.2U W=20U
MP23  21   0  22 100   P12L5   L=1.2U W=20U
MN21  21   0   0   0   N10L5   L=1.0U W=5U
MN22  21  11   0   0   N10L5   L=1.0U W=5U
MN23  21   0   0   0   N10L5   L=1.0U W=5U

MP31  31  21 100 100   P12L5   L=1.2U W=10U
MP32  31 100 100 100   P12L5   L=1.2U W=10U
MN31  31  21  32   0   N10L5   L=1.0U W=5U
MN32  32 100   0   0   N10L5   L=1.0U W=5U

MP41  41  31 100 100   P12L5   L=1.2U W=10U
MN41  41  31   0   0   N10L5   L=1.0U W=5U

C11   11   0  1P
C21   21   0  1P
C31   31   0  1P
C41   41   0  1P
.ENDS

VDD 100    0  5
VIN  1    0  DC 0 PWL(0 0 2N 5)

.TRAN 0.5N 150N
.PRINT TRAN V(1) V(2) V(3) V(4) V(5)
.PRINT TRAN V(11) V(12) V(13) V(41) V(42) V(43)

*.OPTIONS ACCT

**** LEVEL 1 NMOS ****
.MODEL N10L1 NMOS
+ LEVEL=1 TPG=1
+ KP=2.33082E-05
+ LAMBDA=0.013333 VT0=0.69486 GAMMA=0.60309 PHI=1
+ TOX=1.9800000E-08  XJ=0.2U            LD=0.1U           NSUB=4.9999999E+16
+ NSS=0.0000000E+00
+ CJ=4.091E-4        MJ=0.307           PB=1.0
+ CJSW=3.078E-10     MJSW=1.0E-2        
+ CGSO=3.93E-10      CGDO=3.93E-10
**** LEVEL 1 PMOS ****
.MODEL P12L1 PMOS
+ LEVEL=1 TPG=-1
+ KP=7.69968E-06
+ LAMBDA=0.018966 VT0=-0.60865 GAMMA=0.89213 PHI=1
+ TOX=1.9800000E-08  XJ=0.4U            LD=0.28U           NSUB=4.9999999E+17
+ NSS=0.0000000E+00
+ CJ=6.852E-4        MJ=0.429           PB=1.0
+ CJSW=5.217E-10     MJSW=0.351
+ CGSO=7.29E-10      CGDO=7.29E-10
**** LEVEL 3 NMOS ****
.MODEL  N10L3  NMOS
+ LEVEL=3            TPG=+1
+ GAMMA=1.140501     THETA=0.8109787    KAPPA=0.1579183    ETA=5.0622310E-02
+ DELTA=0.000000E+00 UO=812.5126        VMAX=1186662.      VTO=0.8
+ TOX=1.9800000E-08  XJ=0.2U            LD=0.1U            NSUB=4.9999999E+16
+ NSS=0.0000000E+00
+ CJ=4.091E-4        MJ=0.307           PB=1.0
+ CJSW=3.078E-10     MJSW=1.0E-2        
+ CGSO=3.93E-10      CGDO=3.93E-10
**** LEVEL 3 PMOS ****
.MODEL  P12L3  PMOS
+ LEVEL=3            TPG=-1
+ GAMMA=1.211640     THETA=0.1184638    KAPPA=0.2162577    ETA=2.7580135E-02
+ DELTA=0.000000E+00 UO=89.16160        VMAX=5.9000000E+07 VTO=-0.8
+ TOX=1.9800000E-08  XJ=0.4U            LD=0.28U           NSUB=4.9999999E+17
+ NSS=0.0000000E+00
+ CJ=6.852E-4        MJ=0.429           PB=1.0
+ CJSW=5.217E-10     MJSW=0.351
+ CGSO=7.29E-10      CGDO=7.29E-10
**** LEVEL 6 NMOS ****
.MODEL N10L5 NMOS
+ LEVEL=6 TPG=1
+ KC=3.8921e-05 NC=1.1739 KV=0.91602 NV=0.87225
+ LAMBDA0=0.013333 LAMBDA1=0.0046901 VT0=0.69486 GAMMA=0.60309 PHI=1
+ TOX=1.9800000E-08  XJ=0.2U            LD=0.1U           NSUB=4.9999999E+16
+ NSS=0.0000000E+00
+ CJ=4.091E-4        MJ=0.307           PB=1.0
+ CJSW=3.078E-10     MJSW=1.0E-2        
+ CGSO=3.93E-10      CGDO=3.93E-10
**** LEVEL 6 PMOS ****
.MODEL P12L5 PMOS
+ LEVEL=6 TPG=-1
+ KC=6.42696E-06 NC=1.6536 KV=0.92145 NV=0.88345
+ LAMBDA0=0.018966 LAMBDA1=0.0084012 VT0=-0.60865 GAMMA=0.89213 PHI=1
+ TOX=1.9800000E-08  XJ=0.4U            LD=0.28U           NSUB=4.9999999E+17
+ NSS=0.0000000E+00
+ CJ=6.852E-4        MJ=0.429           PB=1.0
+ CJSW=5.217E-10     MJSW=0.351
+ CGSO=7.29E-10      CGDO=7.29E-10
.END
