* simple voltage regulator, example for traditional feedback loop analysis using L and C

Mout out pgate vdd vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=100
R1 out fb 33.3K
R2 fb vss 66.7K

Mp1 mir mir vdd vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=2
Mp2 pgate mir vdd vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=2

M1 pgate set tail vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=10
M2 mir fbinj tail vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=10
Cc pgate vdd 10p

Mb1 tail bn vss vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=4
Mb0 bn bn vss vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=4
Ib vss bn 1u

* breaking the loop with huge inductor
Lloop fb fbinj 100e6
* injecting AC trough huge capacitor
Cinj inj fbinj 100e6
Vinj inj 0 DC 0 AC 1
* load replication for node 'fb' (approximate)
M2rep mirrep fb tailrep vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=10
Mp1rep mirrep mirrep vdd vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=2
Mb1rep tailrep bn vss vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=2


Vset set vss DC 1.2
Vvdd vdd vss DC 3.3
Vvss vss 0 DC 0

Cload out vss 100p
Iload out vss DC 10e-3 PWL 1n 10e-3 2n 1e-3

.model n1 nmos level=49 version=3.3.0 tox=3.5n nch=2.4e17 nsub=5e16 vth0=0.6
.model p1 pmos level=49 version=3.3.0 tox=3.5n nch=2.5e17 nsub=5e16 vth0=-0.7

.option gmin=1e-14 reltol=1e-5 abstol=1e-14
.ac dec 10 1 10e9

.control
ac dec 10 1 10e9
plot db(fb)
.endc
