CMOS 2-STAGE OPERATIONAL AMPLIFIER

VDD 1 0  2.5V
VSS 2 0 -2.5V

IBIAS 9 0 100UA

VPL 3 0 0.0V AC 0.5V
VMI 4 0 0.0V AC 0.5V 180

M1  6 3 5 5 M_PMOS_1 W=15U  L=1U
M2  7 4 5 5 M_PMOS_1 W=15U  L=1U
M3  6 6 2 2 M_NMOS_1 W=7.5U L=1U
M4  7 6 2 2 M_NMOS_1 W=7.5U L=1U
M5  8 7 2 2 M_NMOS_1 W=15U  L=1U
M6  9 9 1 1 M_PMOS_1 W=15U  L=1U
M7  5 9 1 1 M_PMOS_1 W=15U  L=1U
M8  8 9 1 1 M_PMOS_1 W=15U  L=1U

*CC  7 8 0.1PF

.INCLUDE BICMOS.LIB

*.OP
*.AC DEC 10 1K 100G
.DC VPL -5MV 5MV 0.1MV

.OPTIONS ACCT BYPASS=1 METHOD=GEAR
.END
