** NMOSFET: Benchmarking of B4SOI Stress Effect by Jane Xi 05/09/2003.

.option post nopage brief
.option ingold=1
.option gmin=0

m1 d g s 0 p n1 w=1u l=0.1u soimod=0 NF=2 
+SA=0.31u SB=0.2u SD=0.1u 

vg g 0          1.2
vd d 0          1.2 
vs s 0 		0.0
vp p 0 		0.0

.dc vd 0 1.2 0.02 vg 0.4 1.2 0.1 
.include ./nmos4p0.mod
.print dc i(vd)
.end

