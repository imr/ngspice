STATIC LATCH
***   IC=1MA, RE6=3K
***   SPICE ORIGINAL 1-7-80, CIDER REVISED 4-16-93

***   BIAS CIRCUIT
***   RESISTORS
RCC2 6 8 3.33K
REE2 9 0 200
***   TRANSISTORS
Q1 6 8 4 M_NPN1D AREA=8
Q2 8 4 9 M_NPN1D AREA=8

***   MODELS
.INCLUDE BICMOS.LIB

***   SOURCES
VCC 6 0 5V
VREF 3 0 2.5V
VRSET 1 0 PULSE(2V 3V 0.1NS 0.1NS 0.1NS 0.9NS 4NS)
VSET  7 0 PULSE(2V 3V 2.1NS 0.1NS 0.1NS 0.9NS 4NS)

***   LATCH
X1 1 2 3 4 5 6 ECLNOR2
X2 5 7 3 4 2 6 ECLNOR2

***   SUBCIRCUITS
.SUBCKT ECLNOR2 1 2 3 4 5 6
**  RESISTORS
RS 6 11 520
RC2 11 10 900
RE4 12 0 200
RE6 5 0 6K
**  TRANSISTORS
Q1 9 1 8 M_NPN1D AREA=8
Q2 9 2 8 M_NPN1D AREA=8
Q3 11 3 8 M_NPN1D AREA=8
Q4 8 4 12 M_NPN1D AREA=8
Q5 10 10 9 M_NPN1D AREA=8
Q6 6 9 5 M_NPN1D AREA=8
.ENDS ECLNOR2

***   CONTROL CARDS
.TRAN 0.01NS 8NS
.PRINT TRAN V(1) V(7) V(5) V(2)
.OPTIONS ACCT BYPASS=1
.END
