** One-Shot Trigger (Tran): Benchmarking Implementation of BSIM4.7.0 by Mohan V. Dunga 12/13/2006.

Md1 4 in Vdd Vdd  P1 W=3.6u L=0.2u rgeomod=1
Md2 4 in 0 0 N1 W=1.8u L=0.2u rgeomod=1
c4 4 0 100f
Md3 A 4 Vdd Vdd  P1 W=3.6u L=0.2u rgeomod=1 
Md4 A 4 0 0 N1 W=1.8u L=0.2u rgeomod=1
ca a 0 100f

M1 Anot A Vdd Vdd  P1 W=3.6u L=0.2u rgeomod=1
M2 Anot A 0 0 N1 W=1.8u L=0.2u rgeomod=1

M3 Bnot in Vdd Vdd  P1 W=3.6u L=0.2u rgeomod=1
M4 Bnot in 0 0 N1 W=1.8u L=0.2u rgeomod=1

M5 AorBnot 0 Vdd Vdd P1 W=1.8u L=3.6u rgeomod=1
M6 AorBnot in 1 0 N1 W=1.8u L=0.2u rgeomod=1
M7 1 Anot 0 0 N1 W=1.8u L=0.2u

M8 Lnot 0 Vdd Vdd P1 W=1.8u L=3.6u rgeomod=1
M9 Lnot Bnot 2 0 N1 W=1.8u L=0.2u rgeomod=1
M10 2 A 0 0 N1 W=1.8u L=0.2u

M11 out 0 Vdd Vdd P1 W=3.6u L=3.6u rgeomod=1
M12 out AorBnot 3 0 N1 W=1.8u L=0.2u rgeomod=1
M13 3 Lnot 0 0 N1 W=1.8u L=0.2u

Vcc vdd 0 1.8
vin in 0 pulse 0 1.8 1ns .1ns .1ns .8ns 5ns

.include modelcard.nmos
.include modelcard.pmos

.tran 1ns 10ns
.print tran in out
.option post reltol=1e-2 noacct

.end
