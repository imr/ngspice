RC filter
v1 1 0 0 ac 1.0
r1 1 2 1k
c1 2 0 10p
.options noacct
.pz 1 0 2 0 vol pz
.print pz all
.end
