A simple resistor with a voltage source

R1 1 0 10k
V1 1 0 DC 1

.options noacct
.TRAN 1ns 6ns
.PRINT TRAN I(V1)

.END
