Emitter Coupled Pair

VCC	1  0  5v
VEE	2  0  0v
RCP	1  11 10k
RCN	1  21 10k
VBBP	12 0  3v AC 1
VBBN	22 0  3v
IEE	13 2  0.1mA
Q1	11 12 13 M_NPN AREA=8
Q2	21 22 13 M_NPN AREA=8


.MODEL M_NPN nbjt level=2
+ title TWO-DIMENSIONAL NUMERICAL POLYSILICON EMITTER BIPOLAR TRANSISTOR
+ * Since, we are only simulating half of a device, we double the unit width
+ * 1.0 um emitter length
+ options defw=2.0u
+ 
+ *x.mesh w=2.5 n=5
+ x.mesh w=2.0  h.e=0.05 h.m=0.2 r=1.5
+ x.mesh w=0.5  h.s=0.05 h.m=0.1 r=1.5
+ 
+ y.mesh l=-0.2 n=1
+ y.mesh l= 0.0 n=5
+ y.mesh w=0.10 h.e=0.002 h.m=0.01  r=1.5
+ y.mesh w=0.15 h.s=0.002 h.m=0.01  r=1.5
+ y.mesh w=0.35 h.s=0.01  h.m=0.2   r=1.5
+ y.mesh w=0.40 h.e=0.05  h.m=0.2   r=1.5
+ y.mesh w=0.30 h.s=0.05  h.m=0.1   r=1.5
+
+ domain num=1 material=1 x.l=2.0 y.h=0.0
+ domain num=2 material=2 x.h=2.0 y.h=0.0
+ domain num=3 material=3 y.l=0.0
+ material num=1 polysilicon
+ material num=2 oxide
+ material num=3 silicon
+
+ elec num=1 x.l=0.0  x.h=0.0  y.l=1.1  y.h=1.3
+ elec num=2 x.l=0.0  x.h=0.5  y.l=0.0  y.h=0.0
+ elec num=3 x.l=2.0  x.h=3.0  y.l=-0.2 y.h=-0.2
+
+ doping gauss n.type conc=3e20 x.l=2.0 x.h=3.0 y.l=-0.2 y.h=0.0
+ + char.l=0.047 lat.rotate
+ doping gauss p.type conc=1e19 x.l=0.0 x.h=5.0 y.l=-0.2 y.h=0.0
+ + char.l=0.094 lat.rotate
+ doping unif  n.type conc=1e16 x.l=0.0 x.h=5.0 y.l=0.0 y.h=1.3
+ doping gauss n.type conc=5e19 x.l=0.0 x.h=5.0 y.l=1.3 y.h=1.3
+ + char.l=0.100 lat.rotate
+
+ method ac=direct itlim=10
+ models bgn srh auger conctau concmob fieldmob

.OPTIONS ACCT BYPASS=1
.DC VBBP 2.75v 3.25001v 10mv
.PRINT DC V(21) V(11)
.END
