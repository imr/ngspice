VDMOS output

m1 d g s n1
*.model n1 vdmos rb=0.05 is=10n kp=2 bv=12 rd=0.1
.model  N1  vdmos vto=1 cgdmin=0.05p cgdmax=0.2p a=1.2 cgs=0.15p rg=10 kp=2e-4 rb=1e4 is=1e-9 bv=12 cjo=1p ksubthres=0.1

vd d 0 1
vg g 0 1
vs s 0 0

.control
dc vd -2 15 0.05 vg 0 5 1
plot vs#branch
dc vg 0 5 0.05 vd 0.5 2.5 0.5
plot vs#branch ylog
.endc

.end
