test for regression of already fixed bugs

* (exec-spice "ngspice -b %s")

* Bug Tracker
*   #294 B source failure when using an unary minus

b1001_t  n1001_t 0  V=(- (5))
v1001_g  n1001_g 0  -5

v1002_aux aux1002 0 DC=3

b1002_t  n1002_t 0  V=(-(v(aux1002)))
v1002_g  n1002_g 0  -3

.param aux1003=-2

b1003_t  n1003_t 0  V='aux1003**2'
v1003_g  n1003_g 0  4

b1004_t  n1004_t 0  V='-aux1003**2'
v1004_g  n1004_g 0  -4

* unary '+'

b1005_t  n1005_t 0  V=(+ (5))
v1005_g  n1005_g 0  5

b1006_t  n1006_t 0  V=(+(v(aux1002)))
v1006_g  n1006_g 0  3

b1007_t  n1007_t 0  V=+-(5)
v1007_g  n1007_g 0  -5

b1008_t  n1008_t 0  V=-+(5)
v1008_g  n1008_g 0  -5

* ----------------------------------------

.control

define mismatch(a,b,err) abs(a-b)>err

op

let total_count = 0
let fail_count = 0

let tests = 1001 + vector(8)

foreach n $&tests
  set n_test = "n{$n}_t"
  set n_gold = "n{$n}_g"
  if mismatch(v($n_test), v($n_gold), 1e-9)
    let v_test = v($n_test)
    let v_gold = v($n_gold)
    echo "ERROR, test failure, v($n_test) = $&v_test but should be $&v_gold"
    let fail_count = fail_count + 1
  end
  let total_count = total_count + 1
end

if fail_count > 0
  echo "ERROR: $&fail_count of $&total_count tests failed"
  quit 1
else
  echo "INFO: $&fail_count of $&total_count tests failed"
  quit 0
end

.endc

.end
