Multistage filter
v1 1 0 0 ac 1.0
r1 1 2 1k
c1 2 0 10p
e2 3 0 2 0 10
r2 3 4 1k
c2 4 0 1.25p
e3 5 0 4 0 10
r3 5 6 1k
c3 6 0 .02p
.pz 1 0 6 0 vol pz
.print pz all
.end
