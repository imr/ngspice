MOTOROLA MECL III ECL GATE
*.DC VIN -2.0 0 0.02
.TRAN 0.2NS 20NS
VEE 22 0 -6.0
VIN 1 0 PULSE -0.8 -1.8 0.2NS 0.2NS 0.2NS 10NS 20NS
RS 1 2 50
Q1 4 2 6 QMOD AREA = 100P
Q2 4 3 6 QMOD AREA = 100P
Q3 5 7 6 QMOD AREA = 100P
Q4 0 8 7 QMOD AREA = 100P

D1 8 9 DMOD
D2 9 10 DMOD

RP1 3 22 50K
RC1 0 4 100
RC2 0 5 112
RE 6 22 380
R1 7 22 2K
R2 0 8 350
R3 10 22 1958

Q5 0 5 11 QMOD AREA = 100P
Q6 0 4 12 QMOD AREA = 100P

RP2 11 22 560
RP3 12 22 560

Q7 13 12 15 QMOD AREA = 100P
Q8 14 16 15 QMOD AREA = 100P

RE2 15 22 380
RC3 0 13 100
RC4 0 14 112

Q9 0 17 16 QMOD AREA = 100P

R4 16 22 2K
R5 0 17 350
D3 17 18 DMOD
D4 18 19 DMOD
R6 19 22 1958

Q10 0 14 20 QMOD AREA = 100P
Q11 0 13 21 QMOD AREA = 100P

RP4 20 22 560
RP5 21 22 560

.MODEL DMOD D RS=40 TT=0.1NS CJO=0.9PF N=1 IS=1E-14 EG=1.11 VJ=0.8 M=0.5

.MODEL QMOD NBJT LEVEL=1
+ X.MESH NODE=1  LOC=0.0
+ X.MESH NODE=10 LOC=0.9
+ X.MESH NODE=20 LOC=1.1
+ X.MESH NODE=30 LOC=1.4
+ X.MESH NODE=40 LOC=1.6
+ X.MESH NODE=61 LOC=3.0
+ REGION NUM=1 MATERIAL=1
+ MATERIAL NUM=1 SILICON NBGNN=1E17 NBGNP=1E17
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+ DOPING UNIF N.TYPE CONC=1E17 X.L=0.0 X.H=1.0
+ DOPING UNIF P.TYPE CONC=1E16 X.L=0.0 X.H=1.5
+ DOPING UNIF N.TYPE CONC=1E15 X.L=0.0 X.H=3.0
+ MODELS BGNW SRH CONCTAU AUGER CONCMOB FIELDMOB
+ OPTIONS BASE.LENGTH=1.0 BASE.DEPTH=1.25

.OPTIONS ACCT BYPASS=1
.PRINT TRAN V(12) V(21)
.END
