* simple voltage regulator example

Mout out pgate vdd vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=100
R1 out fb 33.3K
R2 fb vss 66.7K

Mp1 mir mir vdd vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=2
Mp2 pgate mir vdd vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=2

M1 pgate set tail vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=10
M2 mir fbinj tail vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=10

Mb1 tail bn vss vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=4
Mb0 bn bn vss vss n1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p m=4
Ib vss bn 1u

Vloop fb fbinj DC 0

Vset set vss DC 1.2 AC 1
Vvdd vdd vss DC 3.3
Vvss vss 0 DC 0

Iload out vss DC 10e-3 PWL 1n 10e-3 2n 9e-3

.model n1 nmos level=49 version=3.3.0 tox=3.5n nch=2.4e17 nsub=5e16 vth0=0.6
.model p1 pmos level=49 version=3.3.0 tox=3.5n nch=2.5e17 nsub=5e16 vth0=-0.7


.loop M2/Gate DEC 10 1 10e9 insrc="Vset" outpos="out" outneg="vss" dir=-1 refnode="set"
.ac dec 10 1 1e9
.tran 1n 10u
