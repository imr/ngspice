Colpitt's Oscillator Circuit
* Colpitt is an harmonic oscillator (LC based) which use
* a capacitive partition of resonator to feed the single 
* active device.
* Predicted frequency is about 3.30435e+06 Hz.

* Models:
.model qnl npn(level=1 bf=80 rb=100 ccs=2pf tf=0.3ns tr=6ns cje=3pf cjc=2pf va=50)

r1 	1 0 	1
q1 	2 1 3	qnl
vcc 	4 0 	5
rl 	4 2 	750
c1 	2 3 	500p
c2 	4 3 	4500p
l1 	4 2 	5uH
re 	3 6 	4.65k
vee 	6 0 	dc -10 pwl 0 0 1e-9 -10 

.control
** transient sim
tran 3n 120u 20u
plot V(2) v(3)
** fft of tran sim
linearize v(3)
fft v(3)
let dbv3 = db(v(3))
plot dbv3 xlimit 1Meg 5Meg
** measure the frequency of oscillation
meas sp fosc MAX_AT dbv3 from=1Meg to=5Meg
** periodic steady state sim
pss 1e6 50e-6 3 256 10 50 5e-3
set xbrushwidth=3
plot v(3) ylimit 0 0.3
.endc

.end




