RTL INVERTER

VIN 1 0 DC 1 PWL 0 4 1NS 0
VCC 12 0 DC 5.0
RC1 12 3 2.5K
RB1 1 2 8K
Q1 3 2 0 QMOD AREA = 100P

.OPTION ACCT BYPASS=1
.TRAN 0.5N 5N
.PRINT TRAN V(2) V(3)

.MODEL QMOD NBJT LEVEL=1
+ X.MESH NODE=1  LOC=0.0
+ X.MESH NODE=61 LOC=3.0
+ REGION NUM=1 MATERIAL=1
+ MATERIAL NUM=1 SILICON NBGNN=1E17 NBGNP=1E17
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+ DOPING UNIF N.TYPE CONC=1E17 X.L=0.0 X.H=1.0
+ DOPING UNIF P.TYPE CONC=1E16 X.L=0.0 X.H=1.5
+ DOPING UNIF N.TYPE CONC=1E15 X.L=0.0 X.H=3.0
+ MODELS BGNW SRH CONCTAU AUGER CONCMOB FIELDMOB
+ OPTIONS BASE.LENGTH=1.0 BASE.DEPTH=1.25

.END
