************  Multiconductor 6-line with ECL drivers  *******
vemm mm g DC -0.4
vepp pp g DC 0.4
vein_left  lin  g PULSE (-0.4 0.4 0N 1N 1N 7N 200N)
vein_right ring g PULSE (-0.4 0.4 2N 1N 1N 7N 200N)

* upper 2 lines
x1 lin g 1 1outn  ECL
x2 mm g 2 2outn   ECL
x7 7 g 7r 7routn  ECL
x8 8 g 8r 8routn  ECL

c7r 7r g 0.1P
c8r 8r g 0.1P

* lower 2 lines
x11 pp g 11 11outn  ECL
x12 rin g 12 12outn  ECL
x5  5 g 5l 5loutn  ECL
x6  6 g 6l 6loutn ECL

c5l 5l g 0.1P
c6l 6l g 0.1P

p1 6 1 2 3 4 5 6   7 8 9 10 11 12 pline
  
.model pline cpl
+C = 0.907067P  -0.657947P -0.0767356P -0.0536544P -0.0386514P -0.0523990P
+   -0.657947P  0.138873P -0.607034P -0.0597635P -0.0258851P -0.0273442P
+   -0.0767356P -0.607034P  1.39328P -0.625675P -0.0425551P -0.0319791P
+   -0.0536544P -0.0597635P -0.625675P  1.07821P -0.255048P -0.0715824P
+   -0.0386514P -0.0258851P -0.0425551P -0.255048P  1.06882P -0.692091P
+   -0.0523990P -0.0273442P -0.0319791P -0.0715824P -0.692091P 0.903603P       
+L = 0.868493E-7 0.781712E-7 0.748428E-7 0.728358E-7 0.700915E-7 0.692178E-7
+    0.781712E-7 0.866074E-7 0.780613E-7 0.748122E-7 0.711591E-7 0.701023E-7
+    0.748428E-7 0.780613E-7 0.865789E-7 0.781095E-7 0.725431E-7 0.711986E-7
+    0.728358E-7 0.748122E-7 0.781095E-7 0.867480E-7 0.744242E-7 0.725826E-7
+    0.700915E-7 0.711591E-7 0.725431E-7 0.744242E-7 0.868022E-7 0.782377E-7
+    0.692178E-7 0.701023E-7 0.711986E-7 0.725826E-7 0.782377E-7 0.868437E-7    
+R = 0.2 0.2 0.2 0.2 0.2 0.2
+G = 0  0  0  0  0  0 
+
+length = 2

*XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX                     
.SUBCKT ECL EIN GND 9 8
*    Input-GND-OUTP-OUTN
RIN  1 2   0.077K
REF  5 6   0.077K
R1   7 N   1.0K
R2   P 3   0.4K
R3   P 4   0.4555K
R4   8 N   0.615K
R5   9 N   0.615K
RL1  8 GND 0.093K
RL2  9 GND 0.093
LIN  EIN 1 0.01U
LREF 5 GND 0.01U
CIN  1 GND 0.68P
CL1  8 GND 1P
CL2  9 GND 1P
Q1 2 3 7 JCNTRAN
Q2 6 4 7 JCNTRAN
Q3 3 P 8 JCNTRAN
Q4 4 P 9 JCNTRAN
VEP  P GND DC 1.25
VEN  N GND DC -3
.ENDS ECL

*.MODEL JCNTRAN (B-C-E)
*XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX                     
.TRAN 0.1N 20N                                               
.PRINT TRAN V(3) V(5) V(8) V(11) V(12)
.MODEL JCNTRAN NPN BF=150 VAF=20V IS=4E-17 RB=300 RC=100 CJE=30FF CJC=30FF
+               CJS=40FF VJE=0.6V VJC=0.6V VJS=0.6 MJE=0.5 MJC=0.5
+               MJS=0.5 TF=16PS TR=1NS
.END
