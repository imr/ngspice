* Capa variable sur la base de la thèse de Marc KODRNJA

.SUBCKT capa 4 6 5 7 8 0
Vref1	26 0	DC 3
Vref2	16 0	DC 3
Vdp	7 0	DC 7
I0	3 0	DC 0.07
Ia1	15 0	DC 0.01
Ia2	25 0	DC 0.01
Ib1	14 0	DC 0.01
Ib2	24 0	DC 0.01

.INCLUDE PN2222.mod
Qv1	4 16 14	PN2222
Qv2	4 26 24	PN2222
Q1	11 14 3	PN2222
Q2	21 24 3	PN2222
Qp1	5 8 11	PN2222
Qm1	6 7 11	PN2222
Qp2	6 8 21	PN2222
Qm2	5 7 21	PN2222
Qc1	4 5 15	PN2222
Qc2	4 6 25	PN2222

R1	4 5	100
R2	4 6	100
C1	15 14	10n
C2	25 24	10n
.ENDS

