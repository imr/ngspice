VBIC Test
VC 1  0 DC 2.0
VB 2  0 DC 0.7
VE 3  0 DC 0.0
*VS 4  0 DC 0.0
Q1 1  2  3  VBIC_HSPICE
.OPTIONS GMIN=1e-13
*.OP
.DC VB 0.2 1.0 0.01

.control
run
plot abs(-i(vc)) abs(-i(vb)) ylimit 1e-12 0.1 ylog
plot abs(-i(vc))/abs(-i(vb)) vs abs(-i(vc)) xlimit 1e-09 0.1 xlog
.endc

.MODEL VBIC NPN LEVEL=4
+ RCX=10 RCI=10 RBX=1 RBI=10 RE=1 RBP=10 RS=10
+ IBEN=1.0E-13
+ RTH=100

.MODEL VBIC_HSPICE NPN LEVEL=4
+ AFN=1 AJC=-0.5 AJE=0.5 AJS=0.5 
+ AVC1=0 AVC2=0 BFN=1 CBCO=0 CBEO=0 CJC=2E-14 
+ CJCP=4E-13 CJE=1E-13 CJEP=1E-13 CTH=0 
+ EA=1.12 EAIC=1.12 EAIE=1.12 EAIS=1.12 EANC=1.12 
+ EANE=1.12 EANS=1.12 FC=0.9 GAMM=2E-11 HRCF=2 
+ IBCI=2E-17 IBCIP=0 IBCN=5E-15 IBCNP=0 
+ IBEI=1E-18 IBEIP=0 IBEN=5E-15 IBENP=0 
+ IKF=2E-3 IKP=2E-4 IKR=2E-4 IS=1E-16 ISP=1E-15 ITF=8E-2 
+ KFN=0 MC=0.33 ME=0.33 MS=0.33 
+ NCI=1 NCIP=1 NCN=2 NCNP=2 NEI=1 NEN=2 
+ NF=1 NFP=1 NR=1 PC=0.75 PE=0.75 PS=0.75 QCO=1E-12 QTF=0 
+ RBI=4 RBP=4 RBX=1 RCI=6 RCX=1 RE=0.2 RS=2 
+ RTH=300 TAVC=0 TD=2E-11 TF=10E-12 TNF=0 TR=100E-12 
+ TNOM=25 VEF=10 VER=4 VO=2 
+ VTF=0 WBE=1 WSP=1 
+ XII=3 XIN=3 XIS=3 XRBI=1 XRCI=1 XRE=1 XRS=1 XTF=20 XVO=0 

.MODEL VBIC_APLAC NPN LEVEL=4 
+ IS=1e-16 IBEI=1e-18 IBEN=5e-15 IBCI=2e-17 IBCN=5e-15 ISP=1e-15 RCX=10
+ RCI=60 RBX=10 RBI=40 RE=2 RS=20 RBP=40 VEF=10 VER=4 IKF=2e-3 ITF=8e-2
+ XTF=20 IKR=2e-4 IKP=2e-4 CJE=1e-13 CJC=2e-14 CJEP=1e-13 CJCP=4e-13 VO=2
+ GAMM=2e-11 HRCF=2 QCO=1e-12 AVC1=2 AVC2=15 TF=10e-12 TR=100e-12 TD=2e-11 RTH=300

.END
