** NMOSFET: Benchmarking Implementation of BSIM4 by Jane Xi 05/09/2003.

** Circuit Description **
m1 2 1 0 0 n1 L=0.09u W=10.0u rgeoMod=1
vgs 1 0 1.2 
vds 2 0 1.2 

.dc vds 0 1.2 0.02 vgs 0 1.2 0.2

.options Temp=-55.0 noacct

.print dc v(1) i(vds)

.include modelcard.nmos
.end
