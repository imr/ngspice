* test ASRC ac analysis with regard to HERTZ and tc1
* (exec-spice "ngspice %s" t)

* Test the implementation of the ASRC device with regard to HERTZ and tc1
* This circuit is deliberatly designed in such a way as to make
*   the original incorrect implementation of the ASRC model obvious,
*   which incorrectly evaluated the ASRC expression for every frequency
*      to recalculate the operating point of the whole circuit
*    instead of calculating the operating point from the expression
*      when HERTZ=0
*   The diode is deliberatly attached here to expose the difference.
* A second aspect is to check the tc1 parameter of the ASRC

.temp 27.0

v0  1 0  dc = 5 ac = 1

b1  1 2  v = 'i(b1) * 1k * (1 + sqrt(hertz/1kHz))' tc1 = 0.01

c2  2 0  30u
d2  2 0  dplain temp=27.0       $ keep diode at 27.0 for simplicity

.model dplain d()

.control

* default is 1e-12, but our golden solution is derived without
set gmin = 0

set reltol = 1e-15
set vntol  = 1e-15
*set abstol = 1e-15
*set chgtol = 1e-24

let uT = boltz * (273.15 + 27.0) / echarge

* These 'boltz' and 'echarge' are literal copied from src/spicelib/devices/dio
*   and differ slightly from our global visible ones
let uT = 1.3806226e-23 / 1.6021918e-19 * (273.15 + 27.0)

op

let u0 = @v0[dc]
let c2 = @c2[capacitance]
let is = @dplain[is]

let gold_r1_dc = 1k * (1 + ($temp - 27.0) * 0.01)

* golden solution of the operating point
*   uT = kT/e
*   i = is * (e^(u/uT - 1)
*   di/du = is * e^~ * kT/e = (i + is) / uT

let cd = 1m
repeat 6
  let f = cd * gold_r1_dc + uT * log(cd/is + 1) - u0
  let f_hat = gold_r1_dc + uT / (cd/is + 1) / is
  let cd = cd - f/f_hat
  let err = cd/-i(v0) - 1
  echo "iteration: err = $&err"
end

let gold_cd = cd
let gold_gd = (cd + is) / uT
let gold_vd = uT * log(cd/is + 1)

let err_cd = @d2[id]/gold_cd - 1
let err_gd = @d2[gd]/gold_gd - 1
let err_vd = @d2[vd]/gold_vd - 1

* compare golden diode model with ngspice solution
* expect errors of several double floating ULP, roughly 1E-15

echo "INFO: err_cd = $&err_cd"
echo "INFO: err_gd = $&err_gd"
echo "INFO: err_vd = $&err_vd"

* now do the 'ac' analysis

ac dec 100 1 1e6

let s = 2*pi*i * frequency

let gold_r1_ac = op1.gold_r1_dc * (1 + sqrt(frequency/1kHz))
let gold_H = 1 / (1 + gold_r1_ac * (s * op1.c2 + op1.gold_gd))

let err = v(2)/gold_H - 1
let err_H = vecmax(abs(err))

echo "INFO: err_H = $&err_H"

* expect errors of several double floating ULP, roughly 1E-15
plot abs(gold_H) abs(v(2))
plot abs(err)

.endc
