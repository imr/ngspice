COLPITT'S OSCILLATOR CIRCUIT

R1 1 0 1
Q1 2 1 3 QMOD AREA = 100P
VCC 4 0 5 
RL 4 2 750
C1 2 3 500P
C2 4 3 4500P
L1 4 2 5UH
RE 3 6 4.65K
VEE 6 0 DC -15 PWL 0 -15 1E-9 -10 

.TRAN 30N 12U
.PRINT TRAN V(2)

.MODEL QMOD NBJT LEVEL=1
+ X.MESH NODE=1  LOC=0.0
+ X.MESH NODE=61 LOC=3.0
+ REGION NUM=1 MATERIAL=1
+ MATERIAL NUM=1 SILICON NBGNN=1E17 NBGNP=1E17
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+ DOPING UNIF N.TYPE CONC=1E17 X.L=0.0 X.H=1.0
+ DOPING UNIF P.TYPE CONC=1E16 X.L=0.0 X.H=1.5
+ DOPING UNIF N.TYPE CONC=1E15 X.L=0.0 X.H=3.0
+ MODELS BGNW SRH CONCTAU AUGER CONCMOB FIELDMOB
+ OPTIONS BASE.LENGTH=1.0 BASE.DEPTH=1.25

.OPTIONS ACCT BYPASS=1
.END
