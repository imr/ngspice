SOA check for bipolar
* LTSPICE or PSPICE compatability must be enabled to correctly parse the
* model below, for example with "set ngbehavior=psa" in .spiceinit.

Vce c 0 -1
Ib b 0 -1u
Ve e 0 0

Q1 c b e MPSA92

.MODEL MPSA92 PNP(IS=9.53E-14 ISE=8.37E-13 ISC=9.99E-11 XTI=3.00 BF=9.80E1 BR=4.78 IKF=3.49E-2 IKR=1.00 XTB=1.5 VAF=2.60E2 VAR=1.40E2 VJE=3.00E-1 VJC=3.00E-1 RE=1.00E-2 RC=1.00E-2 RB=2.76E1 RBM=6.66E-2 IRB=7.02E-4 CJE=9.54E-11 CJC=4.66E-11 .00 FC=5.00E-1 NF=1.00 NR=1.55 NE=1.49 NC=1.50 MJE=4.26E-1 MJC=7.00E-1 TF=9.52E-10 TR=516.9p ITF=4.12E-1 VTF=9.99E5 XTF=1.03 EG=1.11 VCEO=300 ICRATING=500m MFG=SIEMENS pd_max=0.625 rth0=200 tnom=25)

.option warn=1 maxwarns=2
.temp 50

.control
dc Vce 0 -200 -0.1 Ib 0 80u 8u
plot i(Ve)
.endc

.end
