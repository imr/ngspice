Controlled sources test
.tran 2us 5ms
.probe alli

*VCCS
G1 g1 0 2 0 1.5m
RG g1 0 1

*VCVS
E1 e1 0 2 0 2.5m
Re e1 0 1.3

*CCCS
F1 f1 0 vf 3.33
RF f1 0 1

*CCVS
H1 h1 0 vh 4.44
Rh h1 0 1.67

* source control voltage
v2 2 0 DC 0.0 PWL (0 0.9 2e-3 2 4e-3 0.4)
* source control current
I1 3 0 DC 0.0 PWL (0 0 2e-3 2m 4e-3 -2m) $ <--- control current

vf 33 3 dc 0 $ <--- measure the current
vh 0 33 dc 0 $ <--- measure the current
* load voltage


.control
run
display
set xbrushwidth=2

plot i(vh) i(g1) i(h1) i(e1) i(f1)
.endc
.end