.title KiCad schematic
.include "model-card-hicumL0V1p11_mod.lib"
XQ5 GND Net-_R1-Pad2_ A2 VEE DT hicumL0V1p1_c_sbt
Ra2 A2 VEE 510
Rt1 DT GND 1G
V3 In2 GND dc -1.75 pulse(-1.75 -0.9 0 1n 1n 2.5u 5u)
R2 GND Net-_R2-Pad2_ 220
R3 GND Net-_R3-Pad2_ 575
R1 GND Net-_R1-Pad2_ 220
XQ3 Net-_R2-Pad2_ Net-_R3-Pad2_ Net-_Q1-Pad3_ VEE DT hicumL0V1p1_c_sbt
Ra1 A1 VEE 510
XQ4 GND Net-_R2-Pad2_ A1 VEE DT hicumL0V1p1_c_sbt
R4 Net-_R3-Pad2_ VEE 1.92k
XQ1 Net-_R1-Pad2_ IN1 Net-_Q1-Pad3_ VEE DT hicumL0V1p1_c_sbt
XQ2 Net-_R1-Pad2_ IN2 Net-_Q1-Pad3_ VEE DT hicumL0V1p1_c_sbt
R5 Net-_Q1-Pad3_ VEE 780
V2 IN1 GND dc -1.75 pulse(-1.75 -0.9 0 1n 1n 5u 10u)
V1 VEE GND -5.2
.tran 0.1n 100u
.control
pre_osdi test_osdi_win/HICUML0-2.osdi
run
plot a1 a2+2 in1+4 in2+6
.endc
.end
