*** NDINV * 4

VDD 100    0  5
VIN  1    0  DC 0 PWL(0 0 2N 5)

MN10  11 100  12   0   p12l5   L=1.0U W=5U
MN11  11 100  12   0   N10L5   L=1.0U W=5U
MN12  11 100  12   0   N10L1   L=1.0U W=5U

.TRAN 0.5N 150N
.PRINT TRAN V(1) V(2) V(3) V(4) V(5)
.PRINT TRAN V(11) V(12) V(13) V(41) V(42) V(43)
.OPTIONS ACCT

**** LEVEL 1 NMOS ****
.MODEL N10L1 NMOS
+ LEVEL=1 TPG=1
+ KP=2.33082E-05
+ LAMBDA=0.013333 VT0=0.69486 GAMMA=0.60309 PHI=1
+ TOX=1.9800000E-08           LD=0.1U           NSUB=4.9999999E+16
+ NSS=0.0000000E+00
+ CJ=4.091E-4        MJ=0.307           PB=1.0
+ CJSW=3.078E-10     MJSW=1.0E-2        
+ CGSO=3.93E-10      CGDO=3.93E-10
**** LEVEL 6 NMOS ****
.MODEL N10L5 NMOS
+ LEVEL=6 TPG=1
+ KC=3.8921e-05 NC=1.1739 KV=0.91602 NV=0.87225
+ LAMBDA0=0.013333 LAMBDA1=0.0046901 VT0=0.69486 GAMMA=0.60309 PHI=1
+ TOX=1.9800000E-08             LD=0.1U           NSUB=4.9999999E+16
+ NSS=0.0000000E+00
+ CJ=4.091E-4        MJ=0.307           PB=1.0
+ CJSW=3.078E-10     MJSW=1.0E-2        
+ CGSO=3.93E-10      CGDO=3.93E-10
**** LEVEL 6 PMOS ****
.MODEL P12L5 PMOS
+ LEVEL=6 TPG=-1
+ KC=6.42696E-06 NC=1.6536 KV=0.92145 NV=0.88345
+ LAMBDA0=0.018966 LAMBDA1=0.0084012 VT0=-0.60865 GAMMA=0.89213 PHI=1
+ TOX=1.9800000E-08             LD=0.28U           NSUB=4.9999999E+17
+ NSS=0.0000000E+00
+ CJ=6.852E-4        MJ=0.429           PB=1.0
+ CJSW=5.217E-10     MJSW=0.351
+ CGSO=7.29E-10      CGDO=7.29E-10
.END
