TURNOFF TRANSIENT OF PASS TRANSISTOR

M1 11 2 3 4 MMOD W=20UM
CS 1 0 6.0PF
CL 3 0 6.0PF
R1 3 6 200K
VIN 6 0 DC 0
VDRN 1 11 DC 0
VG 2 0 DC 5 PWL 0 5 0.1N 0 1 0
VB 4 0 DC 0.0

.TRAN 0.05NS 0.2NS 0.0NS 0.05NS
.PRINT TRAN V(1) I(VDRN)
.IC V(1)=0 V(3)=0
.OPTION ACCT BYPASS=1

.MODEL MMOD NUMOS
+ X.MESH L=0.0 N=1
+ X.MESH L=0.6 N=4
+ X.MESH L=0.7 N=5
+ X.MESH L=1.0 N=7
+ X.MESH L=1.2 N=11
+ X.MESH L=3.2 N=21
+ X.MESH L=3.4 N=25
+ X.MESH L=3.7 N=27
+ X.MESH L=3.8 N=28
+ X.MESH L=4.4 N=31
+
+ Y.MESH L=-.05 N=1
+ Y.MESH L=0.0  N=5
+ Y.MESH L=.05  N=9
+ Y.MESH L=0.3  N=14
+ Y.MESH L=2.0  N=19
+
+ REGION NUM=1 MATERIAL=1 Y.L=0.0
+ MATERIAL NUM=1 SILICON
+ MOBILITY MATERIAL=1 CONCMOD=SG FIELDMOD=SG
+
+ REGION NUM=2 MATERIAL=2 Y.H=0.0 X.L=0.7 X.H=3.7
+ MATERIAL NUM=2 OXIDE
+
+ ELEC NUM=1 X.L=3.8 X.H=4.4	Y.L=0.0 Y.H=0.0
+ ELEC NUM=2 X.L=0.7 X.H=3.7	IY.L=1  IY.H=1
+ ELEC NUM=3 X.L=0.0 X.H=0.6	Y.L=0.0 Y.H=0.0
+ ELEC NUM=4 X.L=0.0 X.H=4.4	Y.L=2.0 Y.H=2.0
+
+ DOPING UNIF P.TYPE CONC=2.5E16 X.L=0.0 X.H=4.4  Y.L=0.0 Y.H=2.0
+ DOPING UNIF P.TYPE CONC=1E16   X.L=0.0 X.H=4.4  Y.L=0.0 Y.H=0.05
+ DOPING UNIF N.TYPE CONC=1E20   X.L=0.0 X.H=1.1  Y.L=0.0 Y.H=0.2
+ DOPING UNIF N.TYPE CONC=1E20   X.L=3.3 X.H=4.4  Y.L=0.0 Y.H=0.2
+
+ MODELS CONCMOB FIELDMOB
+ METHOD AC=DIRECT ONEC

.END
