* AD22057N SPICE Macro-model         
* Description: Amplifier
* Generic Desc: Bipolar, CSAmp, G=20, BiDir, Auto
* Developed by: ARG / ADSC
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (11/1995)
* Copyright 1995, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
* This version of the AD22057 model simulates the worst-case
* parameters of the 'N' grade. The worst-case parameters
* used correspond to those in the data sheet.
*
* END Notes
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  A1 out
*                |  |  |  |  |  A2 in
*                |  |  |  |  |  |  offset
*                |  |  |  |  |  |  |  output
*                |  |  |  |  |  |  |  |
.SUBCKT AD22057N 1  2  99 50 30 31 40 49
*
* A1 INPUT ATTENUATORS, GAIN, AND OFFSET RESISTORS
*
R1 1 3 200K
R2 2 4 200K
RS1 3 16 1K
RS2 4 18 1K
R3 3 5 41K
R4 4 6 41K
R5 5 6 2.55919K TC=-600U
R6 5 50 250
R7 6 50 250
R8 5 19 9K
R9 6 7 10K
R10 19 40 2K
R11 19 50 2K
R12 7 30 100K
R16 7 50 10K
C1 16 50 5P
C2 17 50 5P
*
* A1 INPUT STAGE AND POLE AT 1MHZ
*
I1 99 8 7.55U
Q1 11 16 9 QP 1
Q2 12 17 10 QP 1
R21 11 50 6.89671K
R22 12 50 6.89671K
R23 8 9 .335
R24 8 10 .335
C3 11 12 11.5P
EOS 61 17 POLY(1) 33 0 -61.149U 1.2
ETC 18 61 POLY(1) 60 0 -49.665M 1
ITC 0 60 49.665U
RTC 60 0 1E3 TC=-107U
*
* GAIN STAGE AND DOMINANT POLE AT 400HZ
*
EREF 98 50 POLY(2) 99 0 50 0 0 0.5 0.5
G1 98 13 12 11 144.997U
R25 13 98 6.89671E6
C4 13 98 57.6923P
D1 13 99 DX
D2 50 13 DX
*
* COMMON MODE STAGE WITH ZERO AT 1KHZ
*
ECM 32 0 POLY(2) 1 0 2 0 0 0.5 0.5
R28 32 33 1E6
R29 33 0 10
CCM 32 33 159P
*
* NEGATIVE ZERO AT 0.6MHZ
*
E1 23 98 13 98 1E6
R26 23 24 1E3
R27 24 98 1E-3
FNZ 23 24 VNZ -1
ENZ 25 98 23 24 1
VNZ 26 98 DC 0
CNZ 25 26 265P
*
* POLE AT 5MHZ
*
G2 98 20 24 98 1E-6
R30 20 98 1E6
C5 20 98 32F
*
* A1 OUTPUT STAGE
*
EIN1 99 27 POLY(1) 20 98 1.5072 1.124
Q216 50 27 28 QP375 3.444
Q218 7 29 99 QP350 9.913
R31 28 29 27K
I2 99 29 4.75U
*
* A2 INPUT STAGE
*
I3 99 34 2.516667U
Q3 35 31 37 QP 1
Q4 36 39 38 QP 1
R32 35 50 106.103K
R33 36 50 106.103K
R34 34 37 85.414K
R35 34 38 85.414K
R13 40 41 20K
R14 41 50 20K
R15 41 49 10K
R17 39 41 95K
*
* A2 1ST GAIN STAGE AND SLEW RATE
*
G3 98 42 36 35 30.159U
R36 42 98 1E6
E2 99 43 POLY(1) 99 98 -0.473 1
E3 44 50 POLY(1) 98 50 -0.473 1
D3 42 43 DX
D4 44 42 DX
*
* A2 2ND GAIN STAGE AND DOMINANT POLE AT 12HZ
*
G4 98 45 42 98 2.5U
R37 45 98 132.629E6
C7 45 98 100P
D5 45 59 DX
D6 55 45 DX
VC1 59 99 5
VC2 50 55 5
*
* NEGATIVE ZERO AT 1MHZ
*
E4 51 98 45 98 1E6
R38 51 52 1E6
R39 52 98 1
FNZ2 51 52 VNZ2 -1
ENZ2 53 98 51 52 1
VNZ2 54 98 0
CNZ2 53 54 159F
*
* A2 OUTPUT STAGE
*
ISY 99 50 469U
EIN2 99 56 POLY(1) 52 98 1.6901 112.132E-3
RIN 46 56 10K
Q316 50 46 47 QP375 1.778
Q310 50 47 48 QP375 5.925
Q318 49 48 57 50 QP350 9.913
I4 99 47 4.75U
I5 99 48 9.5U
VSC 99 57 0
FSC 58 99 VSC 1
QSC 46 58 99 QP350 1
RSC 99 58 89
*
* MODELS USED
*
.MODEL QP350 PNP(IS=1.4E-15 BF=70 CJE=.012P CJC=.06P RE=20 RB=350
+RC=200)
.MODEL QP375 PNP(IS=1.4E-15 CJE=.01P CJC=.05P RE=20 RC=400 RB=100)
.MODEL QP AKO:QP350 PNP(BF=150 VA=100)
.MODEL DX D(CJO=1F RS=.1)
.ENDS

.MODEL QP351 PNP(IS=1.4E-15 BF=70 CJE=.012P CJC=.06P RE=20 RB=350
+RC=200)



