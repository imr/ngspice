** PMOSFET: Benchmarking Implementation of BSIM4.6.1 by Mohan V. Dunga 12/13/2006.

** Circuit Description **
m1 2 1 0 3 p1 L=0.09u W=10.0u rgeoMod=1
vgs 1 0 -1.2
vds 2 0 -0.1
vbs 3 0 0.0

.option noacct
.dc vgs 0.6 -1.2 -0.02 vds -0.1 -1.2 -0.3

.print dc v(2) i(vds)

.include modelcard.pmos 
.end
