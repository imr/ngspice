* pll circuit using xspice code models: version with analog-only iplot
* output frequency 400 MHz
* locked to a 1 or 10 MHz reference

.include shared-pll-xspice.cir

.control
save cont s1 s2 u1n d1 v.xlf.vdd#branch; to save memory
iplot -d 4000 cont
tran 0.1n $&simtime uic
rusage
plot cont s1 s2+1.2 u1n+2.4 d1+3.6 xlimit 4u 5u
plot v.xlf.vdd#branch xlimit 4u 5u ylimit -8m 2m
.endc
.end
