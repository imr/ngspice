EMITTER COUPLED PAIR WITH ACTIVE LOAD

VCC	1 0 5V
VEE	2 0 0V
VINP	4 0 2.99925V  AC 0.5V
VINM	7 0 3V        AC 0.5V 180
IEE	5 2 0.1MA
Q1	3 4 5 M_NPNS AREA=8
Q2	6 7 5 M_NPNS AREA=8
Q3	3 3 1 M_PNPS AREA=8
Q4	6 3 1 M_PNPS AREA=8

.AC DEC 10 10K 100G
.PLOT AC VDB(6)

.INCLUDE BICMOS.LIB

.OPTIONS ACCT RELTOL=1E-6
.END
