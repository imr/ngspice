test if conditions

* test behaviour in special circumstances

v1  1 0  dc 42
R1  1 0  1k


.control

echo "expect Error: missing if condition"
* does not enter cp_istrue()
if
  echo "FAIL: you should not see this"
else
  echo "nonetheless evaluated as FALSE"
end
echo

set testvar_b=""
echo "expect |false|"
* in cp_istrue(): wl!=NULL names==NULL v==NULL
if $testvar_b
  echo "FAIL: you should not see this"
else
  echo "|false|"
end
echo

set testvar_c
echo "expect testvar_c=|TRUE|"
* in cp_istrue(): wl!=NULL names!=NULL v!=NULL
if $testvar_c
  echo "testvar_c=|$testvar_c|"
end
echo

echo "expect Error: testvar_d: no such variable."
echo "expect Warning: NULL arithmetic expression"
* in cp_istrue(): wl!=NULL then wl==NULL names==NULL v==NULL
if $testvar_d
  echo "FAIL: you should not see this"
else
  echo "nonetheless evaluated as FALSE"
end
echo

echo "expect Error(parse.c--checkvalid): testvar_e: no such vector."
* in cp_istrue(): wl!=NULL names==NULL v==NULL
if testvar_e = 3.3
  echo "FAIL: you should not see this"
else
  echo "nonetheless evaluated as FALSE"
end
echo

let testvar_f = 3.5

echo "expect |false|"
if testvar_f = 3.3
  echo "FAIL: you should not see this"
else
  echo "|false|"
end
echo

echo "expect |true|"
if testvar_f = 3.5
  echo "|true|"
else
  echo "FAIL: you should not see this"
end
echo

op
print v(1)

.endc
.end
